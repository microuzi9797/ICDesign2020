`timescale 1ns / 1ps
`define CYCLE 9.1
`define PATTERN 1000

module tb();

//clk generation
reg clk = 1;
always #(`CYCLE/2) clk = ~clk;

//dump waveform
initial begin
	$fsdbDumpfile("sqrt.fsdb");
	$fsdbDumpvars;
end

//time out
initial begin
	#(100000*`CYCLE);
	$display("Simulation time out!");
	$finish;
end

//instatiate DUT
reg rst_n = 1;
reg [9:0] radicand;
wire finish;
wire [4:0] root;
wire [50:0] number;

sqrt DUT(
	.clk(clk),
	.rst_n(rst_n),
	.i_radicand(radicand),
	.o_finish(finish),
	.o_root(root),
	.number(number)
);

//Initial memory
reg [9:0] INPUT_MEM [0:`PATTERN-1];
reg [4:0] GOLDEN_MEM [0:`PATTERN-1];
initial begin
	$readmemb("pattern/radicand.dat", INPUT_MEM);
	$readmemb("pattern/root.dat", GOLDEN_MEM);
end

//Latency
integer latency = 0;
always @(posedge clk or negedge rst_n) begin
	if (~rst_n) begin
		latency = 0;
	end
	else begin
		latency = latency + 1;
	end
end

//input pattern & check result
integer i;
integer err_num = 0;
integer total_latency = 0;

`ifdef PIPELINE
//input
initial begin
	//reset
	@(posedge clk) rst_n = 0;
	@(posedge clk);
	rst_n = 1;
	for (i=0; i<`PATTERN; i=i+1) begin
		#(0.6); //filp flop hold time
		radicand = INPUT_MEM[i];
		@(posedge clk);
	end
end

//check output
integer j;
initial begin
	wait (finish);
	@(negedge clk);
	for (j=0; j<`PATTERN; j=j+1) begin
		if (GOLDEN_MEM[j] === root) begin
			`ifdef DEBUG
				$display("\033[1;92mPattern %3d passed. Input: %4d / Output: %2d / Golden: %2d\033[0m", j, INPUT_MEM[j], root, GOLDEN_MEM[j]);
			`endif
		end
		else begin
			`ifdef DEBUG
				$display("\033[1;31mPattern %3d failed. Input: %4d / Output: %2d / Golden: %2d\033[0m", j, INPUT_MEM[j], root, GOLDEN_MEM[j]);
			`endif
			err_num = err_num + 1;
		end
		@(negedge clk);
	end
	total_latency = latency - 1;

	if (err_num != 0) begin
		USA2;
		$display("\n\033[1;31m=============================================");
		$display("              Simulation failed              ");
		$display("=============================================\033[0m");
	end
	else begin
		USA1;
		$display("\n\033[1;92m=============================================");
		$display("              Simulation passed              ");
		$display("=============================================\033[0m");
	end

	$display("\n\033[1;96m=============================================");
	$display("                   Summary                   ");
	$display("=============================================");
	$display("  	Clock cycle:           %.1f ns", `CYCLE);
	$display("  	Number of transistors: %.0f", $itor(number));
	$display("  	Total excution cycle:  %.0f", $itor(total_latency));
	$display("  	Correctness Score:     %.1f", 40.0 * $itor($itor(`PATTERN) - $itor(err_num)) / $itor(`PATTERN));
	$display("  	Performance Score:     %.1f", $itor(total_latency) * $itor(number) * `CYCLE);
	$display("=============================================\033[0m");

	$finish;
end

`else
initial begin
	for (i=0; i<`PATTERN; i=i+1) begin
		//reset
		@(posedge clk) rst_n = 0;
		@(posedge clk);
		rst_n = 1;
		#(0.6); //filp flop hold time
		radicand = INPUT_MEM[i];

		wait (finish);
		@(negedge clk);
		total_latency = total_latency + latency;
		if (GOLDEN_MEM[i] === root) begin
			`ifdef DEBUG
				$display("\033[1;92mPattern %3d passed. Input: %4d / Output: %2d / Golden: %2d\033[0m", i, INPUT_MEM[i], root, GOLDEN_MEM[i]);
			`endif
		end
		else begin
			`ifdef DEBUG
				$display("\033[1;31mPattern %3d failed. Input: %4d / Output: %2d / Golden: %2d\033[0m", i, INPUT_MEM[i], root, GOLDEN_MEM[i]);
			`endif
			err_num = err_num + 1;
		end
	end

	if (err_num != 0) begin
		BIBLETHUMP;
		$display("\n\033[1;31m=============================================");
		$display("              Simulation failed              ");
		$display("=============================================\033[0m");
	end
	else begin
		POG;
		$display("\n\033[1;92m=============================================");
		$display("              Simulation passed              ");
		$display("=============================================\033[0m");
	end

	$display("\n\033[1;96m=============================================");
	$display("                   Summary                   ");
	$display("=============================================");
	$display("  	Clock cycle:           %.1f ns", `CYCLE);
	$display("  	Number of transistors: %.0f", $itor(number));
	$display("  	Total excution cycle:  %.0f", $itor(total_latency));
	$display("  	Correctness Score:     %.1f", 40.0 * $itor($itor(`PATTERN) - $itor(err_num)) / $itor(`PATTERN));
	$display("  	Performance Score:     %.1f", $itor(total_latency) * $itor(number) * `CYCLE);
	$display("=============================================\033[0m");

	$finish;
end
`endif

task BIBLETHUMP;
begin
	$display("\033[107;40m\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;016m \033[38;5;m&\033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;m#\033[38;5;m#\033[38;5;m/\033[38;5;m,\033[38;5;236m.\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;235m.\033[38;5;236m.\033[38;5;239m*\033[38;5;m/\033[38;5;m#\033[38;5;m%%\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m \033[38;5;m&\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m,\033[38;5;m%%\033[38;5;m(\033[38;5;242m/\033[38;5;236m.\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;236m.\033[38;5;243m/\033[38;5;m#\033[38;5;m&\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m@\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;m(\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;234m \033[38;5;234m \033[38;5;234m \033[38;5;234m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;245m(\033[38;5;m&\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m(\033[38;5;235m.\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;238m,\033[38;5;095m*\033[38;5;138m(\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;181m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;138m(\033[38;5;095m*\033[38;5;238m,\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;236m.\033[38;5;m/\033[38;5;m%%\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;m%%\033[38;5;059m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;095m/\033[38;5;138m(\033[38;5;181m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;175m#\033[38;5;138m#\033[38;5;095m/\033[38;5;238m,\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;240m*\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m&\033[38;5;m/\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;236m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;m*\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m#\033[38;5;239m*\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;095m*\033[38;5;138m(\033[38;5;175m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;175m#\033[38;5;175m#\033[38;5;138m#\033[38;5;095m*\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;m*\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m@\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m%%\033[38;5;240m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;240m*\033[38;5;138m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;095m*\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m,\033[38;5;m%%\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m@\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;138m(\033[38;5;181m%%\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;138m(\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;242m/\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;m@\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m%%\033[38;5;238m,\033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;244m(\033[38;5;181m#\033[38;5;175m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;138m(\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;236m.\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;095m/\033[38;5;175m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;095m/\033[38;5;234m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;m%%\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;138m(\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;239m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;138m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;239m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;m%%\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;246m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;138m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;138m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;m/\033[38;5;m#\033[38;5;m*\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;m#\033[38;5;m@\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;059m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;m(\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;138m(\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;138m(\033[38;5;234m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;245m(\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;138m(\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;138m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;145m#\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m(\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;174m#\033[38;5;138m#\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;138m(\033[38;5;095m/\033[38;5;240m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;240m*\033[38;5;095m/\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;m%%\033[38;5;m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;138m(\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;138m#\033[38;5;095m/\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;138m(\033[38;5;181m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;095m/\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;245m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;095m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;095m/\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m,\033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;238m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;245m(\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;239m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;247m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m/\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;m&\033[38;5;m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;059m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;245m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;m#\033[38;5;m \033[0m");
	$display("\033[38;5;016m \033[38;5;m*\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;138m(\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;243m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;238m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;102m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;m \033[0m");
	$display("\033[38;5;016m \033[38;5;m(\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;244m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;246m(\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;241m*\033[38;5;m,\033[0m");
	$display("\033[38;5;016m \033[38;5;m(\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;238m,\033[38;5;245m(\033[38;5;248m#\033[38;5;102m(\033[38;5;239m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;138m(\033[38;5;240m*\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;095m/\033[38;5;175m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;059m*\033[38;5;m&\033[0m");
	$display("\033[38;5;016m \033[38;5;m(\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;175m#\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m*\033[38;5;234m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;138m(\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;059m*\033[38;5;m/\033[0m");
	$display("\033[38;5;m%%\033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;138m(\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;239m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;138m(\033[38;5;174m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;181m#\033[38;5;138m(\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;240m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;138m(\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;138m(\033[38;5;181m%%\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;138m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;m \033[0m");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;m%%\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m*\033[38;5;181m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;138m#\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m*\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;239m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;095m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;m#\033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;095m/\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;239m*\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;237m,\033[38;5;246m(\033[38;5;174m#\033[38;5;181m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;174m#\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;m&\033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;246m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;095m*\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;067m(\033[38;5;239m,\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;240m*\033[38;5;138m(\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;095m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;138m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;243m/\033[38;5;236m.\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;239m*\033[38;5;073m(\033[38;5;116m#\033[38;5;116m#\033[38;5;109m#\033[38;5;145m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;244m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m/\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;110m#\033[38;5;109m#\033[38;5;109m#\033[38;5;109m#\033[38;5;109m#\033[38;5;109m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;249m#\033[38;5;145m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;138m(\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;237m,\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;145m#\033[38;5;110m#\033[38;5;116m#\033[38;5;110m#\033[38;5;109m#\033[38;5;109m#\033[38;5;073m(\033[38;5;066m(\033[38;5;066m/\033[38;5;066m/\033[38;5;066m(\033[38;5;067m(\033[38;5;109m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m%%\033[38;5;109m#\033[38;5;145m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;234m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;249m#\033[38;5;145m#\033[38;5;175m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;239m,\033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m%%\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;244m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;109m#\033[38;5;116m#\033[38;5;110m#\033[38;5;110m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;110m%%\033[38;5;249m#\033[38;5;175m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m%%\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;145m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;243m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;243m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;242m/\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;110m#\033[38;5;110m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;249m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;181m#\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;m(\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;240m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;109m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;240m*\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;109m#\033[38;5;110m#\033[38;5;249m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;249m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;138m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;145m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;145m#\033[38;5;110m#\033[38;5;109m#\033[38;5;145m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;249m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;138m#\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;m%%\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;095m/\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;249m#\033[38;5;110m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;181m#\033[38;5;145m#\033[38;5;110m#\033[38;5;109m#\033[38;5;145m#\033[38;5;249m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;116m%%\033[38;5;249m%%\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;174m#\033[38;5;138m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;234m.\033[38;5;m#\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m#\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;138m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;145m#\033[38;5;116m%%\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;109m#\033[38;5;109m#\033[38;5;248m#\033[38;5;249m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;109m#\033[38;5;249m%%\033[38;5;174m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;138m(\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;238m,\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m#\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;238m,\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;109m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;145m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;181m#\033[38;5;145m#\033[38;5;109m#\033[38;5;109m#\033[38;5;145m#\033[38;5;249m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;249m#\033[38;5;181m#\033[38;5;181m#\033[38;5;138m#\033[38;5;237m,\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;m#\033[38;5;m&\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m&\033[38;5;241m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;059m*\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;145m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;249m#\033[38;5;109m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;109m#\033[38;5;249m#\033[38;5;138m(\033[38;5;236m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;059m*\033[38;5;m&\033[38;5;m&\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m@\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;237m,\033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;181m#\033[38;5;181m#\033[38;5;145m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;109m#\033[38;5;109m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;110m#\033[38;5;242m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;237m,\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m%%\033[38;5;239m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;238m,\033[38;5;247m#\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;109m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;249m#\033[38;5;109m#\033[38;5;109m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;109m#\033[38;5;237m,\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;238m,\033[38;5;m%%\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;m*\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;066m/\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;249m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;145m#\033[38;5;110m#\033[38;5;109m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;109m#\033[38;5;239m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;247m#\033[38;5;234m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;109m#\033[38;5;110m#\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;116m#\033[38;5;110m#\033[38;5;249m#\033[38;5;145m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;145m#\033[38;5;109m#\033[38;5;249m%%\033[38;5;145m#\033[38;5;145m#\033[38;5;109m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;110m#\033[38;5;116m%%\033[38;5;073m(\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;m#\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;109m#\033[38;5;116m%%\033[38;5;116m#\033[38;5;116m#\033[38;5;116m#\033[38;5;110m#\033[38;5;145m#\033[38;5;145m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;145m#\033[38;5;109m#\033[38;5;110m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;110m#\033[38;5;109m#\033[38;5;066m/\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;242m/\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;241m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;066m/\033[38;5;109m#\033[38;5;116m#\033[38;5;116m#\033[38;5;145m#\033[38;5;145m#\033[38;5;181m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;145m#\033[38;5;249m#\033[38;5;110m%%\033[38;5;249m#\033[38;5;248m#\033[38;5;244m/\033[38;5;236m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;m/\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;244m/\033[38;5;234m.\033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;066m/\033[38;5;109m#\033[38;5;145m#\033[38;5;138m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m#\033[38;5;181m#\033[38;5;247m#\033[38;5;241m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;248m#\033[38;5;m&\033[38;5;m@\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m%%\033[38;5;240m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m \033[38;5;237m,\033[38;5;095m/\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;138m(\033[38;5;095m*\033[38;5;235m.\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;243m/\033[38;5;m%%\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;m%%\033[38;5;m(\033[38;5;236m.\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;240m*\033[38;5;138m(\033[38;5;138m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;175m#\033[38;5;175m#\033[38;5;174m#\033[38;5;138m#\033[38;5;095m/\033[38;5;239m*\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;239m,\033[38;5;m#\033[38;5;m%%\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m \033[38;5;m#\033[38;5;145m#\033[38;5;240m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;238m,\033[38;5;240m*\033[38;5;095m*\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;102m(\033[38;5;102m(\033[38;5;138m(\033[38;5;244m(\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m*\033[38;5;238m,\033[38;5;236m.\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;059m*\033[38;5;m%%\033[38;5;m%%\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m&\033[38;5;m&\033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;m@\033[38;5;m@\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m*\033[38;5;m%%\033[38;5;m(\033[38;5;239m,\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;239m,\033[38;5;m/\033[38;5;m%%\033[38;5;m*\033[38;5;m#\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;m&\033[38;5;m(\033[38;5;m/\033[38;5;m/\033[38;5;m*\033[38;5;236m.\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;235m.\033[38;5;236m.\033[38;5;m,\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m@\033[38;5;m.\033[38;5;m*\033[38;5;m.\033[38;5;m(\033[38;5;m.\033[38;5;m&\033[38;5;m.\033[38;5;m#\033[38;5;m.\033[38;5;m*\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;016m \033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
end
endtask

task UMI;
begin
	$display("\033[107;40m\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;138m(\033[38;5;138m(\033[38;5;241m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;242m/\033[38;5;144m#\033[38;5;180m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;244m(\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;059m*\033[38;5;239m*\033[38;5;059m*\033[38;5;240m*\033[38;5;239m*\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;059m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;243m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;059m*\033[38;5;239m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m#\033[38;5;138m(\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m/\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;242m/\033[38;5;187m&\033[38;5;223m&\033[38;5;180m#\033[38;5;180m#\033[38;5;174m#\033[38;5;138m#\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;138m#\033[38;5;138m#\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;240m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;242m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;240m*\033[38;5;239m,\033[38;5;240m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;241m*\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;244m(\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;247m#\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m/\033[38;5;138m#\033[38;5;095m/\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;241m/\033[38;5;253m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;174m#\033[38;5;138m#\033[38;5;239m*\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;095m/\033[38;5;174m#\033[38;5;138m#\033[38;5;138m(\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;244m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;252m&\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m*\033[38;5;138m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;180m#\033[38;5;180m#\033[38;5;138m#\033[38;5;239m*\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;059m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;240m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;059m*\033[38;5;239m,\033[38;5;239m,\033[38;5;059m*\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;180m#\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;187m&\033[38;5;243m/\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;008m(\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m*\033[38;5;174m#\033[38;5;138m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;243m/\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;144m#\033[38;5;059m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;145m#\033[38;5;180m#\033[38;5;180m#\033[38;5;180m#\033[38;5;138m#\033[38;5;095m/\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;059m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;238m,\033[38;5;242m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;181m%%\033[38;5;144m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;239m*\033[38;5;181m%%\033[38;5;253m&\033[38;5;250m%%\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;138m(\033[38;5;240m*\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;248m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;174m#\033[38;5;144m#\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;249m%%\033[38;5;223m&\033[38;5;181m#\033[38;5;180m#\033[38;5;180m#\033[38;5;174m#\033[38;5;138m(\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;242m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;239m,\033[38;5;238m,\033[38;5;059m*\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;187m&\033[38;5;245m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;180m#\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;251m%%\033[38;5;241m*\033[38;5;239m,\033[38;5;243m/\033[38;5;252m&\033[38;5;187m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;242m/\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;138m#\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;145m#\033[38;5;181m%%\033[38;5;174m#\033[38;5;095m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;243m/\033[38;5;251m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;180m#\033[38;5;138m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;249m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;187m&\033[38;5;180m#\033[38;5;180m#\033[38;5;174m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;060m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;060m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;243m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;252m&\033[38;5;242m/\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;138m(\033[38;5;181m%%\033[38;5;187m&\033[38;5;187m&\033[38;5;252m&\033[38;5;248m#\033[38;5;240m*\033[38;5;239m,\033[38;5;238m,\033[38;5;102m(\033[38;5;252m&\033[38;5;187m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m(\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;251m%%\033[38;5;223m&\033[38;5;180m#\033[38;5;008m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;187m&\033[38;5;253m&\033[38;5;252m&\033[38;5;245m(\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;102m(\033[38;5;251m%%\033[38;5;253m&\033[38;5;187m&\033[38;5;180m#\033[38;5;102m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;250m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;180m%%\033[38;5;180m#\033[38;5;174m#\033[38;5;138m#\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;243m/\033[38;5;095m/\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;095m/\033[38;5;138m#\033[38;5;180m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;252m&\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m/\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;243m/\033[38;5;249m%%\033[38;5;252m&\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;245m(\033[38;5;238m,\033[38;5;238m,\033[38;5;095m/\033[38;5;138m#\033[38;5;101m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;253m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;247m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;253m&\033[38;5;252m&\033[38;5;247m#\033[38;5;241m*\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;180m#\033[38;5;180m#\033[38;5;144m#\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;242m/\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m*\033[38;5;138m(\033[38;5;095m/\033[38;5;101m/\033[38;5;138m(\033[38;5;144m#\033[38;5;181m%%\033[38;5;187m&\033[38;5;253m&\033[38;5;181m&\033[38;5;241m*\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;181m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;181m%%\033[38;5;174m#\033[38;5;095m*\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;247m#\033[38;5;253m&\033[38;5;224m&\033[38;5;187m&\033[38;5;245m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;245m(\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;181m%%\033[38;5;138m(\033[38;5;138m(\033[38;5;181m%%\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;223m&\033[38;5;180m#\033[38;5;180m#\033[38;5;138m#\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;095m/");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;138m#\033[38;5;180m#\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;244m/\033[38;5;238m,\033[38;5;238m,\033[38;5;250m%%\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;187m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;144m#\033[38;5;138m(\033[38;5;138m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;138m(\033[38;5;237m,\033[38;5;238m,\033[38;5;246m(\033[38;5;187m&\033[38;5;144m#\033[38;5;239m*\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;249m#\033[38;5;181m%%\033[38;5;181m%%\033[38;5;181m&\033[38;5;187m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;251m%%\033[38;5;239m,\033[38;5;239m*\033[38;5;250m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;241m*");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;138m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;247m#\033[38;5;238m,\033[38;5;240m*\033[38;5;252m&\033[38;5;249m#\033[38;5;101m/\033[38;5;181m%%\033[38;5;253m&\033[38;5;187m&\033[38;5;187m&\033[38;5;187m&\033[38;5;252m&\033[38;5;252m&\033[38;5;252m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;251m%%\033[38;5;252m&\033[38;5;252m&\033[38;5;253m&\033[38;5;187m&\033[38;5;187m&\033[38;5;187m&\033[38;5;101m/\033[38;5;144m#\033[38;5;102m(\033[38;5;238m,\033[38;5;238m,\033[38;5;252m&\033[38;5;187m&\033[38;5;144m#\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;008m/\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;244m/\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;138m(\033[38;5;144m#\033[38;5;181m&\033[38;5;224m&\033[38;5;223m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;252m&\033[38;5;138m(\033[38;5;138m(\033[38;5;007m%%\033[38;5;239m*\033[38;5;242m/\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;008m(\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;095m/\033[38;5;181m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;144m#\033[38;5;138m(\033[38;5;181m%%\033[38;5;238m,\033[38;5;008m(\033[38;5;181m%%\033[38;5;181m%%\033[38;5;138m(\033[38;5;240m*\033[38;5;235m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;244m(\033[38;5;138m(\033[38;5;138m(\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;246m(\033[38;5;239m,\033[38;5;244m/\033[38;5;253m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;251m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;238m,\033[38;5;239m,\033[38;5;251m%%\033[38;5;187m&\033[38;5;252m&\033[38;5;251m%%\033[38;5;138m(\033[38;5;059m*\033[38;5;236m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m \033[38;5;234m \033[38;5;234m \033[38;5;234m.\033[38;5;234m.\033[38;5;237m,\033[38;5;095m/\033[38;5;145m#\033[38;5;239m,\033[38;5;252m%%\033[38;5;187m&\033[38;5;181m%%\033[38;5;138m(\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;144m#\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;252m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;138m(\033[38;5;181m%%\033[38;5;187m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;102m(\033[38;5;235m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;239m*\033[38;5;244m/\033[38;5;247m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;247m#\033[38;5;248m#\033[38;5;247m#\033[38;5;243m/\033[38;5;234m.\033[38;5;233m \033[38;5;235m.\033[38;5;181m%%\033[38;5;224m&\033[38;5;253m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;252m&\033[38;5;102m(\033[38;5;239m*\033[38;5;249m%%\033[38;5;224m&\033[38;5;253m&\033[38;5;251m%%\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;241m*\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;007m%%\033[38;5;239m,\033[38;5;239m,\033[38;5;008m(\033[38;5;251m%%\033[38;5;236m.\033[38;5;234m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;235m.\033[38;5;238m,\033[38;5;240m*\033[38;5;242m/\033[38;5;059m*\033[38;5;059m*\033[38;5;238m,\033[38;5;236m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;236m.\033[38;5;247m#\033[38;5;187m&\033[38;5;253m&\033[38;5;253m&\033[38;5;144m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;138m(\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;241m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;238m,\033[38;5;251m%%\033[38;5;253m&\033[38;5;187m&\033[38;5;138m(\033[38;5;181m%%\033[38;5;187m&\033[38;5;253m&\033[38;5;252m&\033[38;5;095m/\033[38;5;241m*\033[38;5;234m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;240m*\033[38;5;248m#\033[38;5;145m#\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;248m#\033[38;5;250m%%\033[38;5;243m/\033[38;5;235m.\033[38;5;237m,\033[38;5;251m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;243m/\033[38;5;240m*\033[38;5;253m&\033[38;5;224m&\033[38;5;253m&\033[38;5;248m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;251m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;059m*\033[38;5;239m*\033[38;5;145m#\033[38;5;095m*\033[38;5;249m%%\033[38;5;235m.\033[38;5;240m*\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;246m(\033[38;5;059m*\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;241m*\033[38;5;246m(\033[38;5;248m#\033[38;5;243m/\033[38;5;248m#\033[38;5;245m(\033[38;5;235m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;237m,\033[38;5;007m%%\033[38;5;253m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;145m#\033[38;5;240m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;241m*\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;243m/\033[38;5;187m&\033[38;5;253m&\033[38;5;223m&\033[38;5;253m&\033[38;5;249m#\033[38;5;138m#\033[38;5;251m%%\033[38;5;238m,\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;246m(\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;102m(\033[38;5;248m#\033[38;5;249m%%\033[38;5;249m#\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;095m/\033[38;5;238m,\033[38;5;236m.\033[38;5;233m \033[38;5;235m.\033[38;5;247m(\033[38;5;145m#\033[38;5;249m#\033[38;5;249m#\033[38;5;252m&\033[38;5;224m&\033[38;5;252m&\033[38;5;101m(\033[38;5;144m#\033[38;5;138m#\033[38;5;253m&\033[38;5;224m&\033[38;5;253m&\033[38;5;243m/\033[38;5;242m/\033[38;5;253m&\033[38;5;224m&\033[38;5;253m&\033[38;5;243m/\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;059m*\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;248m#\033[38;5;239m,\033[38;5;102m(\033[38;5;252m&\033[38;5;244m/\033[38;5;145m#\033[38;5;253m&\033[38;5;007m%%\033[38;5;250m%%\033[38;5;007m%%\033[38;5;249m%%\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;253m&\033[38;5;095m/\033[38;5;094m*\033[38;5;058m,\033[38;5;058m,\033[38;5;234m.\033[38;5;234m \033[38;5;008m/\033[38;5;145m#\033[38;5;145m#\033[38;5;248m#\033[38;5;247m#\033[38;5;237m,\033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;235m.\033[38;5;244m/\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;138m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;059m*\033[38;5;242m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;252m%%\033[38;5;223m&\033[38;5;187m&\033[38;5;138m(\033[38;5;187m&\033[38;5;252m&\033[38;5;240m*\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;237m,\033[38;5;247m#\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;248m#\033[38;5;247m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;249m#\033[38;5;094m*\033[38;5;058m,\033[38;5;058m,\033[38;5;237m,\033[38;5;233m \033[38;5;237m,\033[38;5;188m&\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;244m/\033[38;5;247m#\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;239m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;145m#\033[38;5;138m(\033[38;5;224m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;144m#\033[38;5;094m*\033[38;5;094m,\033[38;5;094m,\033[38;5;058m,\033[38;5;058m,\033[38;5;234m.\033[38;5;237m,\033[38;5;248m#\033[38;5;249m%%\033[38;5;145m#\033[38;5;145m#\033[38;5;248m#\033[38;5;237m,\033[38;5;233m \033[38;5;233m \033[38;5;234m.\033[38;5;007m%%\033[38;5;181m%%\033[38;5;181m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;242m/\033[38;5;243m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;059m*\033[38;5;187m&\033[38;5;223m&\033[38;5;187m&\033[38;5;187m&\033[38;5;247m#\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;234m \033[38;5;246m(\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;145m#\033[38;5;007m%%\033[38;5;254m@\033[38;5;251m%%\033[38;5;237m,\033[38;5;251m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;252m&\033[38;5;239m*\033[38;5;234m \033[38;5;233m \033[38;5;236m.\033[38;5;058m,\033[38;5;058m,\033[38;5;237m,\033[38;5;233m \033[38;5;102m(\033[38;5;254m@\033[38;5;255m@\033[38;5;254m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;144m#\033[38;5;248m#\033[38;5;253m&\033[38;5;224m&\033[38;5;251m%%\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;248m#\033[38;5;253m&\033[38;5;224m&\033[38;5;253m&\033[38;5;138m(\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;188m&\033[38;5;255m@\033[38;5;254m@\033[38;5;243m/\033[38;5;236m.\033[38;5;244m(\033[38;5;188m&\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;240m*\033[38;5;235m.\033[38;5;235m.\033[38;5;058m,\033[38;5;094m,\033[38;5;094m,\033[38;5;094m,\033[38;5;058m,\033[38;5;234m \033[38;5;246m(\033[38;5;252m&\033[38;5;249m%%\033[38;5;249m#\033[38;5;249m#\033[38;5;145m#\033[38;5;244m/\033[38;5;233m \033[38;5;233m \033[38;5;234m.\033[38;5;007m%%\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;242m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m/\033[38;5;243m/\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;249m%%\033[38;5;187m&\033[38;5;223m&\033[38;5;187m&\033[38;5;241m*\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;236m,\033[38;5;247m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;251m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;102m(\033[38;5;234m.\033[38;5;238m,\033[38;5;094m,\033[38;5;094m*\033[38;5;094m*\033[38;5;058m,\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;095m/\033[38;5;130m*\033[38;5;094m,\033[38;5;234m.\033[38;5;239m,\033[38;5;254m&\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;144m#\033[38;5;253m&\033[38;5;253m&\033[38;5;243m/\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;243m/\033[38;5;253m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;181m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m@\033[38;5;255m@\033[38;5;254m@\033[38;5;243m/\033[38;5;234m \033[38;5;058m,\033[38;5;094m*\033[38;5;130m/\033[38;5;095m/\033[38;5;234m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;234m \033[38;5;094m*\033[38;5;094m*\033[38;5;094m,\033[38;5;058m,\033[38;5;234m \033[38;5;248m#\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;249m#\033[38;5;145m#\033[38;5;245m(\033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;252m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;247m#\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;243m/\033[38;5;095m/\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;252m&\033[38;5;187m&\033[38;5;187m&\033[38;5;237m,\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;238m,\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;249m#\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;252m%%\033[38;5;234m.\033[38;5;237m,\033[38;5;094m,\033[38;5;130m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;137m/\033[38;5;131m/\033[38;5;137m/\033[38;5;173m(\033[38;5;137m/\033[38;5;137m/\033[38;5;095m/\033[38;5;234m.\033[38;5;102m(\033[38;5;254m@\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;224m&\033[38;5;007m%%\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;252m&\033[38;5;235m.\033[38;5;239m*\033[38;5;131m/\033[38;5;137m/\033[38;5;179m#\033[38;5;137m(\033[38;5;137m/\033[38;5;095m*\033[38;5;131m/\033[38;5;137m(\033[38;5;137m(\033[38;5;131m/\033[38;5;131m/\033[38;5;237m,\033[38;5;236m.\033[38;5;188m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;249m%%\033[38;5;248m#\033[38;5;240m*\033[38;5;233m \033[38;5;233m \033[38;5;239m*\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;248m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;241m*\033[38;5;243m/\033[38;5;101m/\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;187m&\033[38;5;181m%%\033[38;5;239m,\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;236m.\033[38;5;247m#\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;250m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m&\033[38;5;238m,\033[38;5;237m,\033[38;5;131m/\033[38;5;130m/\033[38;5;173m(\033[38;5;179m#\033[38;5;179m#\033[38;5;215m%%\033[38;5;179m#\033[38;5;173m(\033[38;5;222m%%\033[38;5;180m#\033[38;5;235m.\033[38;5;243m/\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;239m*\033[38;5;240m*\033[38;5;252m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;235m.\033[38;5;235m.\033[38;5;137m(\033[38;5;173m#\033[38;5;179m#\033[38;5;179m#\033[38;5;179m#\033[38;5;179m#\033[38;5;180m%%\033[38;5;186m%%\033[38;5;101m/\033[38;5;235m.\033[38;5;243m/\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m&\033[38;5;249m%%\033[38;5;245m(\033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;249m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;145m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;008m/\033[38;5;101m/\033[38;5;101m/\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;237m,\033[38;5;187m%%\033[38;5;144m#\033[38;5;236m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;239m*\033[38;5;248m#\033[38;5;145m#\033[38;5;145m#\033[38;5;250m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;254m&\033[38;5;245m(\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;237m,\033[38;5;235m.\033[38;5;237m,\033[38;5;249m#\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;251m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;188m&\033[38;5;249m%%\033[38;5;239m*\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;240m*\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;102m(\033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;239m,\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;248m#\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;241m*\033[38;5;101m/\033[38;5;101m(\033[38;5;244m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m,\033[38;5;187m&\033[38;5;181m%%\033[38;5;248m#\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;236m,\033[38;5;248m#\033[38;5;248m#\033[38;5;145m#\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;138m(\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m&\033[38;5;059m*\033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;247m#\033[38;5;187m&\033[38;5;224m&\033[38;5;253m&\033[38;5;246m(\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;008m(\033[38;5;101m(\033[38;5;101m(\033[38;5;243m/\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;252m&\033[38;5;187m&\033[38;5;223m&\033[38;5;007m%%\033[38;5;234m.\033[38;5;232m \033[38;5;233m \033[38;5;102m(\033[38;5;248m#\033[38;5;145m#\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;249m%%\033[38;5;235m.\033[38;5;238m,\033[38;5;251m%%\033[38;5;187m&\033[38;5;181m%%\033[38;5;252m&\033[38;5;224m&\033[38;5;187m&\033[38;5;059m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;008m/\033[38;5;244m(\033[38;5;244m(\033[38;5;101m(\033[38;5;059m*\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;251m%%\033[38;5;237m,\033[38;5;234m.\033[38;5;242m/\033[38;5;248m#\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;254m@\033[38;5;248m#\033[38;5;244m(\033[38;5;007m%%\033[38;5;252m&\033[38;5;144m#\033[38;5;095m/\033[38;5;144m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;138m#\033[38;5;248m#\033[38;5;252m&\033[38;5;250m%%\033[38;5;245m(\033[38;5;251m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;247m#\033[38;5;251m%%\033[38;5;224m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;102m(\033[38;5;102m(\033[38;5;102m(\033[38;5;101m/\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;243m/");
	$display("\033[38;5;235m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;252m&\033[38;5;145m#\033[38;5;242m/\033[38;5;252m&\033[38;5;254m&\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;007m%%\033[38;5;247m#\033[38;5;251m%%\033[38;5;224m&\033[38;5;253m&\033[38;5;138m#\033[38;5;181m%%\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;181m%%\033[38;5;253m&\033[38;5;252m&\033[38;5;248m#\033[38;5;249m%%\033[38;5;224m@\033[38;5;224m@\033[38;5;224m@\033[38;5;224m@\033[38;5;224m&\033[38;5;254m&\033[38;5;250m%%\033[38;5;188m&\033[38;5;252m&\033[38;5;138m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;246m(\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;102m(\033[38;5;102m(\033[38;5;102m(\033[38;5;244m(\033[38;5;059m*\033[38;5;238m,\033[38;5;238m,\033[38;5;059m*\033[38;5;102m(");
	$display("\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;224m&\033[38;5;253m&\033[38;5;144m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;144m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;144m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;059m*\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;059m*\033[38;5;102m(\033[38;5;102m(\033[38;5;138m(\033[38;5;102m(\033[38;5;008m(\033[38;5;238m,\033[38;5;239m*\033[38;5;240m*\033[38;5;008m(\033[38;5;138m(");
	$display("\033[38;5;138m(\033[38;5;181m%%\033[38;5;145m#\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;243m/\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;245m(\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;239m*\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;241m/\033[38;5;245m(\033[38;5;245m(\033[38;5;138m(\033[38;5;138m(\033[38;5;102m(\033[38;5;239m,\033[38;5;239m,\033[38;5;059m*\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;237m,\033[38;5;248m#\033[38;5;187m&\033[38;5;251m%%\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;243m/\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;251m%%\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;247m#\033[38;5;244m/\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;243m/\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;102m(\033[38;5;240m*\033[38;5;239m,\033[38;5;243m/\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;237m,\033[38;5;238m,\033[38;5;138m(\033[38;5;138m(\033[38;5;059m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;242m/\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;252m&\033[38;5;247m#\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;242m/\033[38;5;238m,\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;138m#\033[38;5;095m/\033[38;5;237m,\033[38;5;138m(\033[38;5;174m#\033[38;5;138m(\033[38;5;095m/\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;059m*\033[38;5;252m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;239m*\033[38;5;246m(\033[38;5;252m&\033[38;5;249m#\033[38;5;238m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;240m*\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;241m*\033[38;5;239m*\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;137m(\033[38;5;138m#\033[38;5;138m(\033[38;5;237m,\033[38;5;138m(\033[38;5;174m#\033[38;5;137m(\033[38;5;181m%%\033[38;5;243m/\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;252m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;102m(\033[38;5;247m#\033[38;5;250m%%\033[38;5;247m#\033[38;5;245m(\033[38;5;250m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;239m*\033[38;5;102m(\033[38;5;253m&\033[38;5;187m&\033[38;5;247m#\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;238m,\033[38;5;245m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;239m*\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;253m&\033[38;5;187m&\033[38;5;101m/\033[38;5;101m/\033[38;5;240m*\033[38;5;138m(\033[38;5;138m(\033[38;5;187m&\033[38;5;223m&\033[38;5;251m%%\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;251m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;238m,\033[38;5;237m,\033[38;5;240m*\033[38;5;248m#\033[38;5;252m&\033[38;5;188m&\033[38;5;254m@\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;255m@\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;254m@\033[38;5;254m@\033[38;5;254m@\033[38;5;254m@\033[38;5;254m&\033[38;5;253m&\033[38;5;246m(\033[38;5;238m,\033[38;5;237m,\033[38;5;138m(\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;138m(\033[38;5;138m(\033[38;5;224m&\033[38;5;253m&\033[38;5;224m&\033[38;5;245m(\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;008m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;095m/\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;187m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;101m/\033[38;5;144m#\033[38;5;187m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;251m%%\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;247m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;138m(\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;144m#\033[38;5;145m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;241m/\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;245m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;095m/\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;095m/\033[38;5;095m/\033[38;5;138m#\033[38;5;095m/\033[38;5;187m&\033[38;5;253m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;241m*\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;249m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;138m(\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;249m%%\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;008m(\033[38;5;102m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(");
	$display("\033[38;5;187m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;138m(\033[38;5;138m#\033[38;5;095m/\033[38;5;137m(\033[38;5;138m#\033[38;5;187m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m#\033[38;5;095m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;249m%%\033[38;5;241m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;246m(\033[38;5;187m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;138m(\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;252m&\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;246m(\033[38;5;138m(\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;144m#\033[38;5;138m#\033[38;5;138m(\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#\033[38;5;138m#");
	$display("\033[38;5;240m*\033[38;5;252m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;138m#\033[38;5;138m#\033[38;5;138m(\033[38;5;137m/\033[38;5;174m#\033[38;5;138m#\033[38;5;101m/\033[38;5;253m&\033[38;5;223m&\033[38;5;180m#\033[38;5;138m#\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;247m#\033[38;5;251m%%\033[38;5;245m(\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;249m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m,\033[38;5;236m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;145m#\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;252m&\033[38;5;239m*\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;240m*\033[38;5;250m%%\033[38;5;250m%%\033[38;5;138m(\033[38;5;138m#\033[38;5;138m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;138m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;138m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;241m*\033[38;5;181m%%\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;095m/\033[38;5;138m(\033[38;5;174m#\033[38;5;138m(\033[38;5;131m/\033[38;5;138m(\033[38;5;138m#\033[38;5;138m(\033[38;5;223m&\033[38;5;223m&\033[38;5;180m#\033[38;5;174m#\033[38;5;138m(\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;059m*\033[38;5;251m%%\033[38;5;187m&\033[38;5;252m&\033[38;5;138m(\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;247m#\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;095m*\033[38;5;095m*\033[38;5;095m/\033[38;5;095m/\033[38;5;095m/\033[38;5;095m*\033[38;5;095m*\033[38;5;239m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;144m#\033[38;5;239m*\033[38;5;239m*\033[38;5;102m(\033[38;5;252m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;245m(\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m*\033[38;5;250m%%\033[38;5;187m&\033[38;5;187m&\033[38;5;223m&\033[38;5;138m#\033[38;5;137m/\033[38;5;174m#\033[38;5;138m#\033[38;5;095m/\033[38;5;180m#\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;180m#\033[38;5;181m%%\033[38;5;249m%%\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;243m/\033[38;5;252m&\033[38;5;187m&\033[38;5;253m&\033[38;5;187m&\033[38;5;252m&\033[38;5;251m%%\033[38;5;138m(\033[38;5;241m*\033[38;5;239m,\033[38;5;243m/\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;223m&\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m/\033[38;5;239m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;138m(\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;145m#\033[38;5;253m&\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;101m/\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;145m#\033[38;5;187m&\033[38;5;253m&\033[38;5;253m&\033[38;5;181m&\033[38;5;144m#\033[38;5;187m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;180m#\033[38;5;174m#\033[38;5;181m&\033[38;5;223m&\033[38;5;187m&\033[38;5;252m&\033[38;5;138m#\033[38;5;240m*\033[38;5;240m*\033[38;5;250m%%\033[38;5;253m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;187m&\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;174m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;131m(\033[38;5;095m*\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;240m*\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;101m/\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;181m%%\033[38;5;187m&\033[38;5;223m&\033[38;5;187m&\033[38;5;187m&\033[38;5;102m(\033[38;5;240m*\033[38;5;240m*\033[38;5;059m*\033[38;5;144m#\033[38;5;181m&\033[38;5;223m&\033[38;5;187m&\033[38;5;181m&\033[38;5;180m#\033[38;5;181m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;252m&\033[38;5;253m&\033[38;5;138m(\033[38;5;138m#\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;131m(\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;101m/\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;095m/\033[38;5;144m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;253m&\033[38;5;253m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;240m*\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;239m,\033[38;5;187m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;244m/\033[38;5;059m*\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;095m*\033[38;5;138m#\033[38;5;180m#\033[38;5;223m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;095m*\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;248m#\033[38;5;248m#\033[38;5;243m/\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;145m#\033[38;5;240m*\033[38;5;239m*\033[38;5;247m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;138m#\033[38;5;138m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;245m(\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;243m/\033[38;5;145m#\033[38;5;247m#\033[38;5;252m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;247m#\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;247m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;101m/\033[38;5;174m#\033[38;5;180m#\033[38;5;187m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;101m/\033[38;5;251m%%\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;188m&\033[38;5;253m&\033[38;5;250m%%\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;252m&\033[38;5;242m/\033[38;5;240m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m*\033[38;5;242m/\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;138m(\033[38;5;095m/\033[38;5;138m(\033[38;5;174m#\033[38;5;180m#\033[38;5;187m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;138m#\033[38;5;252m&\033[38;5;188m&\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;101m(\033[38;5;254m@\033[38;5;254m&\033[38;5;247m#\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;253m&\033[38;5;246m(\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;095m/\033[38;5;138m(\033[38;5;138m#\033[38;5;180m#\033[38;5;181m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;137m(\033[38;5;253m&\033[38;5;254m&\033[38;5;254m&\033[38;5;138m(\033[38;5;174m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;138m(\033[38;5;254m&\033[38;5;255m@\033[38;5;254m@\033[38;5;245m(\033[38;5;252m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;253m&\033[38;5;252m&\033[38;5;102m(\033[38;5;237m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;102m(\033[38;5;144m#\033[38;5;144m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;137m(\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;138m(\033[38;5;254m&\033[38;5;255m@\033[38;5;254m@\033[38;5;255m@\033[38;5;188m&\033[38;5;145m#\033[38;5;138m(\033[38;5;095m/\033[38;5;131m/\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;138m(\033[38;5;131m(\033[38;5;131m/\033[38;5;244m(\033[38;5;138m#\033[38;5;252m&\033[38;5;188m&\033[38;5;254m@\033[38;5;255m@\033[38;5;254m@\033[38;5;255m@\033[38;5;254m@\033[38;5;145m#\033[38;5;181m%%\033[38;5;253m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;187m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;239m*\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;247m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;239m*\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;137m(\033[38;5;095m/\033[38;5;174m#\033[38;5;144m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;144m#\033[38;5;138m(\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;224m@\033[38;5;224m&\033[38;5;248m#\033[38;5;144m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;144m#\033[38;5;095m/\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;243m/\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;137m(\033[38;5;095m*\033[38;5;138m#\033[38;5;174m#\033[38;5;180m#\033[38;5;181m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m@\033[38;5;224m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;181m%%\033[38;5;217m%%\033[38;5;181m%%\033[38;5;181m%%\033[38;5;217m%%\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;138m#\033[38;5;059m*\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;246m(\033[38;5;144m#\033[38;5;248m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;138m#\033[38;5;095m/\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;224m&\033[38;5;223m&\033[38;5;187m&\033[38;5;181m%%\033[38;5;144m#\033[38;5;138m(\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;138m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m#\033[38;5;138m(\033[38;5;095m*\033[38;5;137m(\033[38;5;174m#\033[38;5;144m#\033[38;5;144m#\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;224m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;181m%%\033[38;5;138m#\033[38;5;138m(\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;095m/\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;137m/\033[38;5;095m*\033[38;5;095m/\033[38;5;138m(\033[38;5;174m#\033[38;5;174m#\033[38;5;180m#\033[38;5;180m%%\033[38;5;181m%%\033[38;5;217m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;180m%%\033[38;5;174m#\033[38;5;138m#\033[38;5;138m(\033[38;5;239m*\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;144m#\033[38;5;248m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#\033[38;5;144m#");
	$display("\033[0");
end
endtask

task POGGERS;
begin
	$display("\033[107;40m\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;m(\033[38;5;243m/\033[38;5;239m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;059m*\033[38;5;244m/\033[38;5;m(\033[38;5;m(\033[38;5;m#\033[38;5;m%%\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m%%\033[38;5;m#\033[38;5;245m(\033[38;5;242m/\033[38;5;240m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m,\033[38;5;236m,\033[38;5;237m,\033[38;5;236m,\033[38;5;236m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;239m*\033[38;5;240m*\033[38;5;244m/\033[38;5;m(\033[38;5;m#\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m(\033[38;5;m&\033[38;5;m#\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m/\033[38;5;m(\033[38;5;m#\033[38;5;m*\033[38;5;235m.\033[38;5;237m,\033[38;5;239m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;m/\033[38;5;m#\033[38;5;m&\033[38;5;m&\033[38;5;m&\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;m&\033[38;5;m&\033[38;5;m(\033[38;5;239m,\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;238m,\033[38;5;236m.\033[38;5;236m.\033[38;5;243m/\033[38;5;m%%\033[38;5;m&\033[38;5;m#\033[38;5;m(\033[38;5;m#\033[38;5;m(\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m#\033[38;5;m#\033[38;5;m*\033[38;5;236m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m \033[38;5;234m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;237m,\033[38;5;234m.\033[38;5;237m,\033[38;5;059m*\033[38;5;240m*\033[38;5;235m.\033[38;5;236m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;237m,\033[38;5;237m,\033[38;5;m/\033[38;5;m&\033[38;5;m/\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m&\033[38;5;m#\033[38;5;m%%\033[38;5;248m#\033[38;5;102m(\033[38;5;241m*\033[38;5;237m,\033[38;5;234m \033[38;5;233m \033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;237m,\033[38;5;237m,\033[38;5;243m/\033[38;5;252m%%\033[38;5;m&\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m&\033[38;5;m&\033[38;5;m%%\033[38;5;102m(\033[38;5;239m,\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;236m.\033[38;5;234m \033[38;5;234m.\033[38;5;237m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;236m.\033[38;5;236m,\033[38;5;243m/\033[38;5;m#\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m&\033[38;5;145m#\033[38;5;240m*\033[38;5;236m.\033[38;5;236m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;237m,\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;236m.\033[38;5;234m.\033[38;5;236m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;235m.\033[38;5;239m*\033[38;5;m#\033[38;5;m&\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m \033[38;5;m&\033[38;5;m%%\033[38;5;240m*\033[38;5;235m.\033[38;5;238m,\033[38;5;239m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;238m,\033[38;5;243m/\033[38;5;247m#\033[38;5;250m%%\033[38;5;252m&\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;252m&\033[38;5;249m#\033[38;5;244m(\033[38;5;240m*\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;236m.\033[38;5;239m,\033[38;5;239m,\033[38;5;235m.\033[38;5;235m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;240m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;238m,\033[38;5;235m.\033[38;5;234m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;237m,\033[38;5;234m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;239m*\033[38;5;m#\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m%%\033[38;5;m%%\033[38;5;238m,\033[38;5;234m.\033[38;5;235m.\033[38;5;238m,\033[38;5;102m(\033[38;5;251m%%\033[38;5;254m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;243m/\033[38;5;236m.\033[38;5;236m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;235m.\033[38;5;234m.\033[38;5;239m,\033[38;5;065m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;239m*\033[38;5;243m/\033[38;5;248m#\033[38;5;252m&\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;253m&\033[38;5;250m%%\033[38;5;245m(\033[38;5;059m*\033[38;5;236m.\033[38;5;236m,\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;237m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;234m.\033[38;5;241m*\033[38;5;m%%\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m&\033[38;5;247m#\033[38;5;240m*\033[38;5;059m*\033[38;5;250m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;252m&\033[38;5;247m#\033[38;5;059m*\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;238m,\033[38;5;242m/\033[38;5;248m#\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;239m,\033[38;5;236m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;237m,\033[38;5;234m \033[38;5;237m,\033[38;5;102m(\033[38;5;252m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;243m/\033[38;5;236m.\033[38;5;236m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;234m.\033[38;5;235m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;236m.\033[38;5;m#\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m&\033[38;5;246m(\033[38;5;239m*\033[38;5;245m(\033[38;5;254m&\033[38;5;255m@\033[38;5;253m&\033[38;5;243m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;236m.\033[38;5;246m(\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;248m#\033[38;5;236m,\033[38;5;236m.\033[38;5;236m,\033[38;5;240m*\033[38;5;145m#\033[38;5;255m@\033[38;5;188m&\033[38;5;247m#\033[38;5;239m,\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;235m.\033[38;5;240m*\033[38;5;247m#\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;244m(\033[38;5;236m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;235m.\033[38;5;236m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;236m.\033[38;5;m(\033[38;5;m&\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m%%\033[38;5;m*\033[38;5;059m*\033[38;5;250m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;239m*\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;238m,\033[38;5;242m/\033[38;5;252m&\033[38;5;254m@\033[38;5;247m#\033[38;5;236m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;237m,\033[38;5;247m#\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;247m#\033[38;5;237m,\033[38;5;237m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;237m,\033[38;5;245m(\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m&\033[38;5;242m/\033[38;5;240m*\033[38;5;250m%%\033[38;5;254m&\033[38;5;255m@\033[38;5;252m&\033[38;5;240m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;243m/\033[38;5;251m%%\033[38;5;188m&\033[38;5;252m&\033[38;5;245m(\033[38;5;234m.\033[38;5;233m \033[38;5;244m(\033[38;5;253m&\033[38;5;251m%%\033[38;5;240m*\033[38;5;232m \033[38;5;233m \033[38;5;243m/\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;243m/\033[38;5;239m,\033[38;5;249m%%\033[38;5;255m@\033[38;5;252m&\033[38;5;059m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;240m*\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;244m(\033[38;5;240m*\033[38;5;239m,\033[38;5;237m,\033[38;5;236m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;237m,\033[38;5;m#\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m&\033[38;5;m@\033[38;5;m@\033[38;5;m%%\033[38;5;240m*\033[38;5;243m/\033[38;5;251m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;252m&\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m,\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;239m*\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;243m/\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;246m(\033[38;5;237m,\033[38;5;249m#\033[38;5;255m@\033[38;5;188m&\033[38;5;243m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;238m,\033[38;5;248m#\033[38;5;253m&\033[38;5;254m@\033[38;5;252m&\033[38;5;102m(\033[38;5;235m.\033[38;5;232m \033[38;5;241m/\033[38;5;253m&\033[38;5;255m@\033[38;5;249m%%\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;243m/\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;252m&\033[38;5;245m(\033[38;5;235m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;241m*\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m&\033[38;5;242m/\033[38;5;240m*\033[38;5;249m%%\033[38;5;188m&\033[38;5;255m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;236m.\033[38;5;239m,\033[38;5;236m,\033[38;5;233m \033[38;5;016m \033[38;5;237m,\033[38;5;102m(\033[38;5;239m*\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;238m,\033[38;5;059m*\033[38;5;188m&\033[38;5;015m@\033[38;5;253m&\033[38;5;241m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;249m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;246m(\033[38;5;234m \033[38;5;232m \033[38;5;234m.\033[38;5;236m.\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;242m/\033[38;5;235m.\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;247m#\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m#\033[38;5;m&\033[38;5;m*\033[38;5;239m*\033[38;5;145m#\033[38;5;254m&\033[38;5;015m@\033[38;5;255m@\033[38;5;252m&\033[38;5;243m/\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;237m,\033[38;5;246m(\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;250m%%\033[38;5;236m.\033[38;5;239m*\033[38;5;252m&\033[38;5;015m@\033[38;5;254m@\033[38;5;246m(\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;243m/\033[38;5;250m%%\033[38;5;251m%%\033[38;5;248m#\033[38;5;241m*\033[38;5;234m \033[38;5;016m \033[38;5;234m \033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;246m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;246m(\033[38;5;241m*\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;236m.\033[38;5;242m/\033[38;5;m&\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m \033[38;5;m&\033[38;5;m&\033[38;5;m%%\033[38;5;m#\033[38;5;240m*\033[38;5;059m*\033[38;5;250m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;102m(\033[38;5;239m*\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;241m*\033[38;5;247m#\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;244m/\033[38;5;237m,\033[38;5;237m,\033[38;5;240m*\033[38;5;235m.\033[38;5;243m/\033[38;5;188m&\033[38;5;015m@\033[38;5;255m@\033[38;5;246m(\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;246m(\033[38;5;246m(\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;246m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;254m@\033[38;5;248m#\033[38;5;239m*\033[38;5;235m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;238m,\033[38;5;007m%%\033[38;5;m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;m@\033[38;5;m#\033[38;5;m&\033[38;5;m&\033[38;5;m(\033[38;5;237m,\033[38;5;239m,\033[38;5;246m(\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;253m&\033[38;5;249m%%\033[38;5;243m/\033[38;5;238m,\033[38;5;235m.\033[38;5;238m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;235m.\033[38;5;239m*\033[38;5;007m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;254m&\033[38;5;247m#\033[38;5;236m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m,\033[38;5;245m(\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;239m*\033[38;5;236m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;235m.\033[38;5;247m#\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;102m(\033[38;5;235m.\033[38;5;238m,\033[38;5;240m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;239m,\033[38;5;059m*\033[38;5;243m/\033[38;5;246m(\033[38;5;249m#\033[38;5;250m%%\033[38;5;251m%%\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;252m&\033[38;5;007m%%\033[38;5;249m%%\033[38;5;247m#\033[38;5;102m(\033[38;5;243m/\033[38;5;240m*\033[38;5;238m,\033[38;5;236m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;236m.\033[38;5;238m,\033[38;5;246m(\033[38;5;188m&\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;252m&\033[38;5;248m#\033[38;5;244m(\033[38;5;241m*\033[38;5;239m*\033[38;5;239m*\033[38;5;241m*\033[38;5;243m/\033[38;5;247m#\033[38;5;251m%%\033[38;5;254m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;248m#\033[38;5;240m*\033[38;5;236m,\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;242m/\033[38;5;m&\033[38;5;m.\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m%%\033[38;5;239m,\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m,\033[38;5;240m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;243m/\033[38;5;007m%%\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;188m&\033[38;5;249m%%\033[38;5;243m/\033[38;5;237m,\033[38;5;236m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;239m*\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m*\033[38;5;m*\033[38;5;m%%\033[38;5;m#\033[38;5;243m/\033[38;5;239m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m,\033[38;5;236m,\033[38;5;236m.\033[38;5;236m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;234m.\033[38;5;237m,\033[38;5;065m/\033[38;5;240m*\033[38;5;238m,\033[38;5;236m.\033[38;5;234m.\033[38;5;236m.\033[38;5;059m*\033[38;5;245m(\033[38;5;250m%%\033[38;5;188m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;251m%%\033[38;5;246m(\033[38;5;241m*\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;236m.\033[38;5;234m.\033[38;5;236m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;236m.\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;m%%\033[38;5;m/\033[38;5;239m*\033[38;5;236m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;235m.\033[38;5;234m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m,\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m%%\033[38;5;m#\033[38;5;241m*\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;238m,\033[38;5;236m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;247m#\033[38;5;237m,\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;240m*\033[38;5;236m.\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;242m/\033[38;5;235m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;239m,\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;102m(\033[38;5;236m.\033[38;5;239m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;235m.\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m#\033[38;5;238m,\033[38;5;237m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;237m,\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;053m,\033[38;5;089m,\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m*\033[38;5;089m,\033[38;5;237m,\033[38;5;236m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;237m,\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;236m.\033[38;5;235m.\033[38;5;m%%\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m(\033[38;5;239m,\033[38;5;236m.\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;236m.\033[38;5;053m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;125m*\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;239m,\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;239m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;236m.\033[38;5;238m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;236m.\033[38;5;236m.\033[38;5;m%%\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m%%\033[38;5;243m/\033[38;5;237m,\033[38;5;239m*\033[38;5;131m*\033[38;5;131m*\033[38;5;239m,\033[38;5;235m.\033[38;5;053m,\033[38;5;161m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;236m.\033[38;5;239m*\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m/\033[38;5;m@\033[38;5;m%%\033[38;5;239m*\033[38;5;238m,\033[38;5;131m*\033[38;5;131m/\033[38;5;095m*\033[38;5;239m,\033[38;5;234m.\033[38;5;089m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;161m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;053m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;238m,\033[38;5;235m.\033[38;5;234m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;m/\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m/\033[38;5;m@\033[38;5;m&\033[38;5;244m(\033[38;5;237m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;235m.\033[38;5;089m*\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;053m,\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;237m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;237m,\033[38;5;234m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;235m.\033[38;5;247m#\033[38;5;m,\033[38;5;m,\033[38;5;m&\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m&\033[38;5;246m(\033[38;5;237m,\033[38;5;239m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;236m.\033[38;5;237m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;053m,\033[38;5;236m.\033[38;5;234m.\033[38;5;236m.\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;236m.\033[38;5;235m.\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;238m,\033[38;5;007m%%\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m*\033[38;5;m&\033[38;5;245m(\033[38;5;237m,\033[38;5;239m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;235m.\033[38;5;237m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;237m,\033[38;5;234m.\033[38;5;238m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;239m*\033[38;5;235m.\033[38;5;236m.\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;236m.\033[38;5;242m/\033[38;5;m%%\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m@\033[38;5;m&\033[38;5;244m(\033[38;5;237m,\033[38;5;239m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;236m.\033[38;5;053m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;236m.\033[38;5;235m.\033[38;5;239m*\033[38;5;131m*\033[38;5;131m*\033[38;5;239m,\033[38;5;234m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;246m(\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m(\033[38;5;m%%\033[38;5;244m/\033[38;5;237m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;236m.\033[38;5;089m,\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;089m,\033[38;5;237m,\033[38;5;234m.\033[38;5;237m,\033[38;5;095m*\033[38;5;131m*\033[38;5;095m*\033[38;5;235m.\033[38;5;235m.\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;236m.\033[38;5;m*\033[38;5;m#\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;243m/\033[38;5;237m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;239m*\033[38;5;235m.\033[38;5;089m*\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;089m,\033[38;5;053m,\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;236m.\033[38;5;239m*\033[38;5;095m*\033[38;5;131m/\033[38;5;095m*\033[38;5;237m,\033[38;5;234m.\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;236m.\033[38;5;247m#\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;241m*\033[38;5;236m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;238m,\033[38;5;236m.\033[38;5;125m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;236m.\033[38;5;234m.\033[38;5;235m.\033[38;5;239m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;236m.\033[38;5;236m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;238m,\033[38;5;235m.\033[38;5;243m/\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;059m*\033[38;5;237m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;236m.\033[38;5;237m,\033[38;5;125m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;053m,\033[38;5;235m.\033[38;5;238m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;236m.\033[38;5;235m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;235m.\033[38;5;242m/\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m#\033[38;5;059m*\033[38;5;239m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;235m.\033[38;5;053m,\033[38;5;161m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m*\033[38;5;089m,\033[38;5;235m.\033[38;5;236m.\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;237m,\033[38;5;235m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;235m.\033[38;5;241m/\033[38;5;m&\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m#\033[38;5;240m*\033[38;5;239m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;239m*\033[38;5;235m.\033[38;5;089m*\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;089m*\033[38;5;236m,\033[38;5;235m.\033[38;5;239m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;236m.\033[38;5;235m.\033[38;5;239m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;235m.\033[38;5;244m(\033[38;5;m&\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;240m*\033[38;5;239m,\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;238m,\033[38;5;236m.\033[38;5;125m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m*\033[38;5;237m,\033[38;5;235m.\033[38;5;237m,\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;235m.\033[38;5;236m.\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;237m,\033[38;5;m%%\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;240m*\033[38;5;238m,\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;238m,\033[38;5;235m.\033[38;5;125m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;167m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;125m/\033[38;5;089m,\033[38;5;235m.\033[38;5;236m.\033[38;5;239m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;238m,\033[38;5;235m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;237m,\033[38;5;237m,\033[38;5;102m(\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;240m*\033[38;5;239m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m*\033[38;5;237m,\033[38;5;236m,\033[38;5;125m*\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;125m/\033[38;5;089m*\033[38;5;236m.\033[38;5;235m.\033[38;5;238m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;236m.\033[38;5;235m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;237m,\033[38;5;236m,\033[38;5;244m/\033[38;5;m&\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;240m*\033[38;5;237m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;237m,\033[38;5;235m.\033[38;5;237m,\033[38;5;125m*\033[38;5;167m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m/\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;125m*\033[38;5;238m,\033[38;5;235m.\033[38;5;235m.\033[38;5;239m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;237m,\033[38;5;234m.\033[38;5;235m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m,\033[38;5;244m(\033[38;5;m%%\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;242m/\033[38;5;237m,\033[38;5;239m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m/\033[38;5;095m*\033[38;5;239m*\033[38;5;237m,\033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;053m,\033[38;5;089m*\033[38;5;125m*\033[38;5;161m/\033[38;5;167m/\033[38;5;167m/\033[38;5;167m/\033[38;5;168m/\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;168m(\033[38;5;167m/\033[38;5;167m/\033[38;5;125m*\033[38;5;089m*\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;239m*\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;235m.\033[38;5;237m,\033[38;5;247m#\033[38;5;m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m#\033[38;5;m*\033[38;5;237m,\033[38;5;239m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;239m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;m/\033[38;5;m#\033[38;5;m.\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m,\033[38;5;m%%\033[38;5;239m*\033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;239m,\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;238m,\033[38;5;236m.\033[38;5;234m.\033[38;5;236m.\033[38;5;238m,\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;059m*\033[38;5;m#\033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m&\033[38;5;m#\033[38;5;238m,\033[38;5;236m.\033[38;5;238m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;095m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m,\033[38;5;235m.\033[38;5;235m.\033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;239m*\033[38;5;239m*\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;237m,\033[38;5;243m/\033[38;5;m#\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m@\033[38;5;m%%\033[38;5;243m/\033[38;5;236m.\033[38;5;236m,\033[38;5;238m,\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;239m,\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;240m*\033[38;5;102m(\033[38;5;145m#\033[38;5;m%%\033[38;5;m&\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m/\033[38;5;m%%\033[38;5;245m(\033[38;5;239m*\033[38;5;236m.\033[38;5;236m,\033[38;5;238m,\033[38;5;239m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;240m*\033[38;5;m/\033[38;5;m(\033[38;5;249m%%\033[38;5;m%%\033[38;5;m*\033[38;5;m/\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;m#\033[38;5;m&\033[38;5;m#\033[38;5;m/\033[38;5;m*\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;239m*\033[38;5;240m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;065m*\033[38;5;240m*\033[38;5;239m*\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;237m,\033[38;5;236m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;239m*\033[38;5;m*\033[38;5;m/\033[38;5;m#\033[38;5;m%%\033[38;5;m%%\033[38;5;m&\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;016m \033[38;5;m.\033[38;5;m.\033[38;5;m&\033[38;5;m \033[38;5;m%%\033[38;5;m&\033[38;5;m&\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m(\033[38;5;247m#\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;246m(\033[38;5;247m#\033[38;5;247m#\033[38;5;m(\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m&\033[38;5;m&\033[38;5;m&\033[38;5;m,\033[38;5;m(\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m#\033[38;5;m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[0m");
end
endtask

task POG;
begin
	$display("\033[107;40m\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;188m&\033[38;5;238m,\033[38;5;236m,\033[38;5;248m#\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;250m%%\033[38;5;243m/\033[38;5;234m.\033[38;5;245m(\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;239m,\033[38;5;236m,\033[38;5;236m.\033[38;5;236m,\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;188m&\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;231m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;233m \033[38;5;238m,\033[38;5;234m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;236m.\033[38;5;237m,\033[38;5;243m/\033[38;5;241m*\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;235m.\033[38;5;254m&\033[38;5;253m&\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;240m*\033[38;5;253m&\033[38;5;239m,\033[38;5;235m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;240m*\033[38;5;237m,\033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;242m/\033[38;5;247m#\033[38;5;236m.\033[38;5;234m.\033[38;5;234m.\033[38;5;236m.\033[38;5;251m%%\033[38;5;255m@\033[38;5;248m#\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;236m,\033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;236m.\033[38;5;240m*\033[38;5;235m.\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;252m&\033[38;5;236m.\033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m \033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m \033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;243m/\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m \033[38;5;234m \033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;252m&\033[38;5;255m@\033[38;5;255m@\033[38;5;145m#\033[38;5;239m*\033[38;5;255m@\033[38;5;242m/\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;238m,\033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;236m.\033[38;5;236m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;252m&\033[38;5;254m@\033[38;5;247m#\033[38;5;243m/\033[38;5;241m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;231m@\033[38;5;251m%%\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;251m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;237m,\033[38;5;239m,\033[38;5;145m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;253m&\033[38;5;239m*\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;052m.\033[38;5;236m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;052m.\033[38;5;052m.\033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;238m,\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;102m(\033[38;5;235m.\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;233m \033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;236m.\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;173m#\033[38;5;173m(\033[38;5;174m#\033[38;5;216m%%\033[38;5;210m#\033[38;5;174m#\033[38;5;173m#\033[38;5;173m(\033[38;5;131m/\033[38;5;095m*\033[38;5;052m,\033[38;5;052m.\033[38;5;052m.\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;244m(\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;243m/\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m*\033[38;5;238m,\033[38;5;094m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;173m#\033[38;5;173m(\033[38;5;131m/\033[38;5;131m*\033[38;5;094m,\033[38;5;052m.\033[38;5;052m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m.\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;239m,\033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;237m,\033[38;5;095m*\033[38;5;131m(\033[38;5;137m(\033[38;5;131m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m#\033[38;5;216m#\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;131m/\033[38;5;094m,\033[38;5;052m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;244m/\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;233m \033[38;5;234m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;235m.\033[38;5;238m,\033[38;5;095m*\033[38;5;173m(\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m#\033[38;5;215m#\033[38;5;215m#\033[38;5;215m#\033[38;5;215m#\033[38;5;215m#\033[38;5;209m#\033[38;5;173m#\033[38;5;131m*\033[38;5;052m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;237m,\033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;095m*\033[38;5;137m(\033[38;5;174m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;215m#\033[38;5;215m#\033[38;5;209m#\033[38;5;173m(\033[38;5;052m,\033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;239m,\033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;235m.\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m*\033[38;5;173m(\033[38;5;174m#\033[38;5;173m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;095m*\033[38;5;233m \033[38;5;232m \033[38;5;234m.\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;059m*\033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;235m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;239m*\033[38;5;239m*\033[38;5;094m,\033[38;5;131m(\033[38;5;209m#\033[38;5;173m#\033[38;5;209m#\033[38;5;209m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;173m(\033[38;5;095m*\033[38;5;233m \033[38;5;233m \033[38;5;243m/\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;237m,\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;233m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;215m#\033[38;5;215m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;180m%%\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m(\033[38;5;174m#\033[38;5;180m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m#\033[38;5;174m#\033[38;5;095m*\033[38;5;233m \033[38;5;059m*\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;251m%%\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;234m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;239m*\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;173m(\033[38;5;131m*\033[38;5;094m*\033[38;5;094m,\033[38;5;001m,\033[38;5;052m,\033[38;5;052m,\033[38;5;052m,\033[38;5;052m,\033[38;5;052m,\033[38;5;001m,\033[38;5;001m,\033[38;5;001m,\033[38;5;095m*\033[38;5;131m/\033[38;5;167m(\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;173m#\033[38;5;131m/\033[38;5;094m,\033[38;5;052m.\033[38;5;234m.\033[38;5;235m.\033[38;5;245m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;235m.\033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;235m.\033[38;5;238m,\033[38;5;131m/\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;167m/\033[38;5;167m(\033[38;5;173m(\033[38;5;174m#\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;173m(\033[38;5;131m/\033[38;5;095m*\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;238m,\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;145m#\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;235m.\033[38;5;239m,\033[38;5;131m/\033[38;5;173m#\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;209m#\033[38;5;209m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;173m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m#\033[38;5;210m#\033[38;5;173m#\033[38;5;138m#\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;095m*\033[38;5;173m(\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;174m#\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;167m(\033[38;5;167m/\033[38;5;167m/\033[38;5;167m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;173m(\033[38;5;167m(\033[38;5;167m/\033[38;5;167m/\033[38;5;173m(\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m#\033[38;5;174m#\033[38;5;255m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;007m%%\033[38;5;234m.\033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;238m,\033[38;5;131m/\033[38;5;174m(\033[38;5;167m(\033[38;5;131m/\033[38;5;239m*\033[38;5;052m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;095m*\033[38;5;173m(\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;209m#\033[38;5;167m/\033[38;5;130m*\033[38;5;131m*\033[38;5;131m(\033[38;5;174m#\033[38;5;180m#\033[38;5;181m%%\033[38;5;101m/\033[38;5;235m.\033[38;5;052m.\033[38;5;052m,\033[38;5;131m*\033[38;5;131m/\033[38;5;167m/\033[38;5;167m(\033[38;5;173m(\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;131m*\033[38;5;052m,\033[38;5;052m.\033[38;5;052m.\033[38;5;238m,\033[38;5;101m/\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m,\033[38;5;173m(\033[38;5;131m/\033[38;5;088m,\033[38;5;124m*\033[38;5;124m*\033[38;5;130m*\033[38;5;131m/\033[38;5;167m(\033[38;5;131m/\033[38;5;001m,\033[38;5;052m.\033[38;5;052m.\033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;234m.\033[38;5;235m.\033[38;5;234m.\033[38;5;236m.\033[38;5;239m*\033[38;5;131m/\033[38;5;137m(\033[38;5;210m#\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;174m#\033[38;5;174m(\033[38;5;052m,\033[38;5;052m.\033[38;5;094m,\033[38;5;094m*\033[38;5;167m(\033[38;5;173m(\033[38;5;216m#\033[38;5;216m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;174m#\033[38;5;167m(\033[38;5;167m(\033[38;5;131m/\033[38;5;210m#\033[38;5;217m%%\033[38;5;217m&\033[38;5;138m(\033[38;5;234m.\033[38;5;236m.\033[38;5;145m#\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;248m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;131m/\033[38;5;210m#\033[38;5;131m*\033[38;5;167m/\033[38;5;210m#\033[38;5;216m%%\033[38;5;210m#\033[38;5;167m/\033[38;5;131m/\033[38;5;130m*\033[38;5;131m/\033[38;5;131m/\033[38;5;094m*\033[38;5;094m*\033[38;5;094m,\033[38;5;052m,\033[38;5;052m.\033[38;5;234m.\033[38;5;234m \033[38;5;234m.\033[38;5;235m.\033[38;5;236m,\033[38;5;238m,\033[38;5;238m,\033[38;5;095m*\033[38;5;137m(\033[38;5;173m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;210m#\033[38;5;216m%%\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;210m#\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;095m/\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;234m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;052m.\033[38;5;173m(\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;167m/\033[38;5;088m,\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;131m/\033[38;5;095m*\033[38;5;052m.\033[38;5;235m.\033[38;5;235m.\033[38;5;237m,\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;131m/\033[38;5;173m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;167m(\033[38;5;167m(\033[38;5;167m/\033[38;5;167m/\033[38;5;167m(\033[38;5;173m(\033[38;5;209m#\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;216m%%\033[38;5;210m#\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;130m*\033[38;5;130m*\033[38;5;131m*\033[38;5;131m/\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;248m#\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;095m*\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;167m(\033[38;5;130m*\033[38;5;124m,\033[38;5;130m*\033[38;5;130m*\033[38;5;167m/\033[38;5;131m/\033[38;5;167m/\033[38;5;173m(\033[38;5;209m#\033[38;5;173m#\033[38;5;131m(\033[38;5;052m,\033[38;5;052m.\033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;238m,\033[38;5;095m*\033[38;5;131m/\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;216m%%\033[38;5;209m#\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;137m(\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;238m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;095m*\033[38;5;216m%%\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;167m/\033[38;5;167m/\033[38;5;167m(\033[38;5;209m#\033[38;5;167m/\033[38;5;167m(\033[38;5;216m%%\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;173m(\033[38;5;095m*\033[38;5;052m.\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;236m,\033[38;5;095m*\033[38;5;131m/\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;180m#\033[38;5;255m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;095m*\033[38;5;210m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;167m(\033[38;5;210m#\033[38;5;216m%%\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;131m*\033[38;5;052m.\033[38;5;236m.\033[38;5;237m,\033[38;5;236m.\033[38;5;236m.\033[38;5;239m,\033[38;5;095m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;173m#\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;238m,\033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;237m,\033[38;5;137m(\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;131m/\033[38;5;094m*\033[38;5;052m,\033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;131m*\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;216m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m#\033[38;5;174m#\033[38;5;254m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m \033[38;5;095m/\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;209m#\033[38;5;173m(\033[38;5;173m(\033[38;5;131m/\033[38;5;094m*\033[38;5;238m,\033[38;5;237m,\033[38;5;235m.\033[38;5;236m.\033[38;5;236m.\033[38;5;052m.\033[38;5;052m,\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;174m#\033[38;5;174m#\033[38;5;174m#\033[38;5;173m#\033[38;5;173m(\033[38;5;173m(\033[38;5;209m(\033[38;5;209m(\033[38;5;173m(\033[38;5;173m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;138m(\033[38;5;231m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;240m*\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;239m,\033[38;5;095m*\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;131m/\033[38;5;167m/\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;239m*\033[38;5;238m,\033[38;5;237m,\033[38;5;236m,\033[38;5;052m,\033[38;5;094m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;173m(\033[38;5;167m/\033[38;5;130m*\033[38;5;088m,\033[38;5;001m,\033[38;5;001m,\033[38;5;088m,\033[38;5;001m,\033[38;5;001m,\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;173m#\033[38;5;173m(\033[38;5;253m&\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;252m&\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;235m.\033[38;5;239m*\033[38;5;239m*\033[38;5;239m,\033[38;5;058m,\033[38;5;058m,\033[38;5;094m*\033[38;5;131m/\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;131m(\033[38;5;131m(\033[38;5;131m/\033[38;5;131m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m%%\033[38;5;216m%%\033[38;5;174m#\033[38;5;131m/\033[38;5;094m*\033[38;5;094m,\033[38;5;094m*\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;137m(\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;234m.\033[38;5;238m,\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;094m*\033[38;5;094m*\033[38;5;095m*\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;209m#\033[38;5;210m#\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;173m(\033[38;5;167m/\033[38;5;167m(\033[38;5;137m(\033[38;5;144m#\033[38;5;231m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;231m@\033[38;5;253m&\033[38;5;235m.\033[38;5;233m \033[38;5;233m \033[38;5;233m \033[38;5;235m.\033[38;5;239m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;137m(\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m#\033[38;5;210m#\033[38;5;210m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m#\033[38;5;216m%%\033[38;5;210m%%\033[38;5;216m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;217m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m%%\033[38;5;210m#\033[38;5;173m(\033[38;5;253m&\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;144m#\033[38;5;095m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;173m(\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;131m(\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;210m#\033[38;5;173m#\033[38;5;167m(\033[38;5;167m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m%%\033[38;5;216m%%\033[38;5;216m%%\033[38;5;174m#\033[38;5;131m/\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;138m(\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;180m#\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;131m*\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;173m(\033[38;5;173m(\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;174m#\033[38;5;210m%%\033[38;5;210m#\033[38;5;174m#\033[38;5;131m/\033[38;5;131m*\033[38;5;052m,\033[38;5;052m.\033[38;5;052m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;052m \033[38;5;052m.\033[38;5;239m,\033[38;5;095m/\033[38;5;101m/\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;137m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;088m*\033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;052m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;233m \033[38;5;234m \033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;095m*\033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;173m(\033[38;5;137m/\033[38;5;137m/\033[38;5;137m(\033[38;5;137m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;167m(\033[38;5;167m(\033[38;5;210m#\033[38;5;210m%%\033[38;5;210m#\033[38;5;131m/\033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;052m.\033[38;5;052m,\033[38;5;001m,\033[38;5;001m,\033[38;5;089m*\033[38;5;095m*\033[38;5;095m/\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;173m(\033[38;5;137m(\033[38;5;137m(\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;173m(\033[38;5;167m/\033[38;5;167m/\033[38;5;167m/\033[38;5;167m(\033[38;5;203m(\033[38;5;203m(\033[38;5;131m/\033[38;5;131m*\033[38;5;088m,\033[38;5;088m,\033[38;5;125m*\033[38;5;124m*\033[38;5;124m*\033[38;5;124m*\033[38;5;131m*\033[38;5;131m/\033[38;5;254m&\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;174m#\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m(\033[38;5;131m/\033[38;5;131m(\033[38;5;131m(\033[38;5;131m(\033[38;5;131m(\033[38;5;137m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;209m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;210m#\033[38;5;209m#\033[38;5;209m#\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m/\033[38;5;167m(\033[38;5;203m(\033[38;5;203m(\033[38;5;204m#\033[38;5;203m#\033[38;5;203m(\033[38;5;203m(\033[38;5;203m(\033[38;5;210m#\033[38;5;167m(\033[38;5;138m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;254m&\033[38;5;174m#\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m#\033[38;5;209m#\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m/\033[38;5;167m(\033[38;5;203m(\033[38;5;203m(\033[38;5;203m(\033[38;5;203m(\033[38;5;173m(\033[38;5;174m#\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;231m@\033[38;5;217m&\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;167m(\033[38;5;167m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;173m(\033[38;5;167m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m*\033[38;5;131m*\033[38;5;095m*\033[38;5;131m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m*\033[38;5;095m/\033[38;5;101m/\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;174m#\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;167m(\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;173m#\033[38;5;173m(\033[38;5;167m(\033[38;5;131m/\033[38;5;095m*\033[38;5;094m*\033[38;5;094m*\033[38;5;094m*\033[38;5;094m*\033[38;5;094m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;137m(\033[38;5;255m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;231m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;224m@\033[38;5;174m#\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;173m(\033[38;5;173m(\033[38;5;173m#\033[38;5;167m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;137m(\033[38;5;254m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;253m&\033[38;5;173m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m/\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m/\033[38;5;131m*\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;138m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;181m%%\033[38;5;174m#\033[38;5;131m(\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;131m/\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;095m*\033[38;5;131m/\033[38;5;137m(\033[38;5;131m/\033[38;5;095m/\033[38;5;138m#\033[38;5;231m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;231m@\033[38;5;255m@\033[38;5;253m&\033[38;5;174m#\033[38;5;174m#\033[38;5;138m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;137m(\033[38;5;131m(\033[38;5;131m(\033[38;5;137m(\033[38;5;138m#\033[38;5;251m%%\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@");
	$display("\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;255m@\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@");
	$display("\033[0");
end
endtask

task USA1;
begin
	$display("\033[107;40m\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;089m*\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;237m,\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;089m*\033[38;5;167m/\033[38;5;131m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;116m&\033[38;5;159m&\033[38;5;067m(\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;116m%%\033[38;5;159m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;116m%%\033[38;5;235m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;234m.\033[38;5;073m#\033[38;5;159m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;123m&\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;058m,\033[38;5;220m#\033[38;5;220m#\033[38;5;094m*\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;003m*\033[38;5;011m%%\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;226m#\033[38;5;058m*\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;234m.\033[38;5;142m/\033[38;5;136m/\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;066m(\033[38;5;159m&\033[38;5;123m&\033[38;5;123m&\033[38;5;159m&\033[38;5;066m/\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;239m*\033[38;5;235m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;242m/\033[38;5;243m/\033[38;5;240m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;116m#\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m#\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;241m*\033[38;5;123m&\033[38;5;123m&\033[38;5;073m#\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;246m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;234m.\033[38;5;073m#\033[38;5;159m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;117m&\033[38;5;234m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;239m*\033[38;5;123m&\033[38;5;123m&\033[38;5;123m&\033[38;5;236m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;246m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;242m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;060m*\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;066m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;116m%%\033[38;5;123m&\033[38;5;159m&\033[38;5;060m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;073m(\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;159m&\033[38;5;067m(\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;184m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;058m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;238m,\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;253m&\033[38;5;224m&\033[38;5;218m&\033[38;5;218m&\033[38;5;181m%%\033[38;5;138m#\033[38;5;242m/\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;246m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;073m(\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m(\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;240m*\033[38;5;155m%%\033[38;5;156m%%\033[38;5;156m%%\033[38;5;192m%%\033[38;5;107m/\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;184m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;132m(\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;224m@\033[38;5;218m&\033[38;5;095m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;239m*\033[38;5;117m%%\033[38;5;117m&\033[38;5;117m&\033[38;5;116m%%\033[38;5;238m,\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;107m/\033[38;5;192m%%\033[38;5;156m%%\033[38;5;149m#\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;058m,\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;136m/\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;181m%%\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;224m@\033[38;5;218m&\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;066m/\033[38;5;123m&\033[38;5;123m&\033[38;5;116m#\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;142m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m(\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;236m.\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;211m%%\033[38;5;138m(\033[38;5;239m*\033[38;5;236m.\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;248m#\033[38;5;102m(\033[38;5;m/\033[38;5;m/\033[38;5;m/\033[38;5;243m/\033[38;5;242m/\033[38;5;239m*\033[38;5;236m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;066m/\033[38;5;159m&\033[38;5;073m#\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;011m%%\033[38;5;178m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;243m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;138m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;238m,\033[38;5;243m/\033[38;5;248m#\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;016m \033[38;5;066m*\033[38;5;073m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;184m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;245m(\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;188m&\033[38;5;015m@\033[38;5;251m%%\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;003m*\033[38;5;011m%%\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;058m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;245m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;016m \033[38;5;016m \033[38;5;243m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;102m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;234m.\033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m(\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;016m \033[38;5;236m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;003m*\033[38;5;011m%%\033[38;5;220m#\033[38;5;220m#\033[38;5;184m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;232m \033[38;5;233m \033[38;5;247m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;142m/\033[38;5;220m#\033[38;5;220m#\033[38;5;226m#\033[38;5;100m*\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;224m@\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;187m%%\033[38;5;217m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;242m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;003m*\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;003m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;237m,\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;234m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;145m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;230m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;095m/\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;089m,\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;138m#\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;234m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;184m(\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;131m/\033[38;5;204m#\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;187m&\033[38;5;237m,\033[38;5;235m.\033[38;5;067m(\033[38;5;232m \033[38;5;233m \033[38;5;181m#\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;136m/\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;235m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;247m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;236m.\033[38;5;234m.\033[38;5;116m%%\033[38;5;066m/\033[38;5;016m \033[38;5;239m,\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;241m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;058m,\033[38;5;220m#\033[38;5;220m#\033[38;5;226m%%\033[38;5;094m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;008m/\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;138m(\033[38;5;016m \033[38;5;239m*\033[38;5;116m&\033[38;5;116m%%\033[38;5;232m \033[38;5;235m.\033[38;5;181m%%\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;233m \033[38;5;016m \033[38;5;233m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;178m(\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;224m@\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;224m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;239m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;244m(\033[38;5;252m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;233m \033[38;5;016m \033[38;5;244m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;016m \033[38;5;235m.\033[38;5;073m#\033[38;5;123m&\033[38;5;123m&\033[38;5;238m,\033[38;5;233m \033[38;5;138m(\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;016m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;058m,\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;224m@\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;247m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m%%\033[38;5;236m.\033[38;5;016m \033[38;5;236m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;181m%%\033[38;5;232m \033[38;5;233m \033[38;5;116m#\033[38;5;123m&\033[38;5;117m&\033[38;5;123m&\033[38;5;059m*\033[38;5;016m \033[38;5;095m/\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;237m,\033[38;5;016m \033[38;5;142m/\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;178m(\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;237m,\033[38;5;149m#\033[38;5;156m%%\033[38;5;234m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;230m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;145m#\033[38;5;234m.\033[38;5;016m \033[38;5;073m#\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;059m*\033[38;5;016m \033[38;5;095m/\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;236m.\033[38;5;232m \033[38;5;136m/\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;003m*\033[38;5;232m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;156m%%\033[38;5;155m%%\033[38;5;149m#\033[38;5;156m%%\033[38;5;149m#\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;224m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;230m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;236m.\033[38;5;232m \033[38;5;116m#\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;236m.\033[38;5;234m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;234m \033[38;5;233m \033[38;5;136m/\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;178m(\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;065m/\033[38;5;192m%%\033[38;5;149m#\033[38;5;149m#\033[38;5;149m#\033[38;5;149m#\033[38;5;192m%%\033[38;5;239m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;239m*\033[38;5;232m \033[38;5;073m(\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m#\033[38;5;016m \033[38;5;237m,\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;233m \033[38;5;232m \033[38;5;136m/\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;184m#\033[38;5;058m,\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;155m%%\033[38;5;156m%%\033[38;5;149m#\033[38;5;149m#\033[38;5;149m#\033[38;5;155m%%\033[38;5;156m%%\033[38;5;239m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;224m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;230m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;016m \033[38;5;239m*\033[38;5;117m%%\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;123m&\033[38;5;237m,\033[38;5;232m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;234m \033[38;5;016m \033[38;5;178m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;136m/\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;107m(\033[38;5;192m%%\033[38;5;155m#\033[38;5;149m#\033[38;5;149m#\033[38;5;149m#\033[38;5;155m%%\033[38;5;192m%%\033[38;5;107m/\033[38;5;m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;234m.\033[38;5;059m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;235m.\033[38;5;234m.\033[38;5;073m#\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m(\033[38;5;232m \033[38;5;235m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;241m*\033[38;5;016m \033[38;5;058m,\033[38;5;226m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;226m%%\033[38;5;142m/\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m,\033[38;5;149m#\033[38;5;192m%%\033[38;5;156m%%\033[38;5;155m#\033[38;5;156m%%\033[38;5;156m%%\033[38;5;192m%%\033[38;5;155m%%\033[38;5;065m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;016m \033[38;5;236m.\033[38;5;116m%%\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;116m%%\033[38;5;235m.\033[38;5;016m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;016m \033[38;5;234m.\033[38;5;142m(\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;058m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;238m,\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;016m \033[38;5;238m,\033[38;5;117m&\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m(\033[38;5;233m \033[38;5;234m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;232m \033[38;5;232m \033[38;5;100m*\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;178m(\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;058m,\033[38;5;149m#\033[38;5;192m%%\033[38;5;192m%%\033[38;5;192m%%\033[38;5;149m#\033[38;5;240m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;243m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;230m@\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;217m&\033[38;5;223m&\033[38;5;217m&\033[38;5;217m&\033[38;5;217m&\033[38;5;223m&\033[38;5;224m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;145m#\033[38;5;016m \033[38;5;238m,\033[38;5;117m&\033[38;5;123m&\033[38;5;117m&\033[38;5;117m&\033[38;5;123m&\033[38;5;073m(\033[38;5;233m \033[38;5;236m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;233m \033[38;5;016m \033[38;5;058m,\033[38;5;226m#\033[38;5;011m%%\033[38;5;136m/\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;101m/\033[38;5;192m%%\033[38;5;156m%%\033[38;5;155m#\033[38;5;192m%%\033[38;5;101m/\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;244m(\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;060m*\033[38;5;123m&\033[38;5;159m&\033[38;5;116m%%\033[38;5;235m.\033[38;5;016m \033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;237m,\033[38;5;192m%%\033[38;5;156m%%\033[38;5;149m#\033[38;5;155m%%\033[38;5;156m%%\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;058m,\033[38;5;156m%%\033[38;5;155m%%\033[38;5;149m#\033[38;5;149m#\033[38;5;192m%%\033[38;5;065m/\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;145m#\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;241m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;149m#\033[38;5;192m%%\033[38;5;149m#\033[38;5;156m%%\033[38;5;107m(\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;233m \033[38;5;100m/\033[38;5;226m%%\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;220m#\033[38;5;235m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;238m,\033[38;5;016m \033[38;5;237m,\033[38;5;138m#\033[38;5;238m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;237m,\033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;246m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;003m*\033[38;5;094m*\033[38;5;058m,\033[38;5;235m.\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;238m,\033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;211m%%\033[38;5;204m#\033[38;5;204m#\033[38;5;131m/\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;252m&\033[38;5;249m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;239m*\033[38;5;016m \033[38;5;234m.\033[38;5;204m#\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;211m%%\033[38;5;204m(\033[38;5;204m(\033[38;5;204m#\033[38;5;204m(\033[38;5;204m(\033[38;5;211m%%\033[38;5;224m@\033[38;5;218m&\033[38;5;138m(\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;234m.\033[38;5;204m#\033[38;5;204m(\033[38;5;205m#\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;211m%%\033[38;5;204m(\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;204m#\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;224m@\033[38;5;096m/\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;145m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;234m.\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;211m#\033[38;5;218m&\033[38;5;218m&\033[38;5;175m%%\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;095m/\033[38;5;181m%%\033[38;5;224m@\033[38;5;095m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;008m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;204m#\033[38;5;204m(\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;236m.\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;243m/\033[38;5;248m#\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;238m,\033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;204m#\033[38;5;204m#\033[38;5;204m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;238m,\033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;204m#\033[38;5;168m(\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;241m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;244m(\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;237m,\033[38;5;016m \033[38;5;237m,\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;204m#\033[38;5;131m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;145m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;236m.\033[38;5;016m \033[38;5;237m,\033[38;5;204m(\033[38;5;211m%%\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;218m&\033[38;5;131m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;240m*\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;244m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;236m.\033[38;5;016m \033[38;5;237m,\033[38;5;204m#\033[38;5;204m(\033[38;5;204m(\033[38;5;211m%%\033[38;5;218m&\033[38;5;218m&\033[38;5;224m&\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;246m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;236m.\033[38;5;016m \033[38;5;237m,\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;204m#\033[38;5;131m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;241m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;059m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;234m.\033[38;5;016m \033[38;5;240m*\033[38;5;224m@\033[38;5;181m%%\033[38;5;236m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;234m.\033[38;5;016m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;242m/\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;241m*\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;016m \033[38;5;233m \033[38;5;247m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;242m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;102m(\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;243m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;145m#\033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;244m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;059m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;243m/\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;240m*\033[38;5;016m \033[38;5;232m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;246m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;246m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;244m/\033[38;5;015m@\033[38;5;252m&\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;252m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;240m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;059m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;239m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;008m(\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;242m/\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m(\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;m@\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[0");
end
endtask

task USA2;
begin
	$display("\033[107;40m\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;239m,\033[38;5;145m#\033[38;5;244m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;234m \033[38;5;102m(\033[38;5;007m%%\033[38;5;059m*\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;242m/\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;102m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m%%\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;239m,\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;239m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;245m(\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;066m/\033[38;5;080m#\033[38;5;073m(\033[38;5;236m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;235m.\033[38;5;080m#\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;245m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;236m.\033[38;5;060m*\033[38;5;237m,\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;246m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;073m(\033[38;5;080m#\033[38;5;023m*\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;244m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;235m.\033[38;5;016m \033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;239m,\033[38;5;238m,\033[38;5;236m.\033[38;5;235m.\033[38;5;233m \033[38;5;233m \033[38;5;236m.\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;073m(\033[38;5;066m/\033[38;5;234m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;237m,\033[38;5;242m/\033[38;5;246m(\033[38;5;007m%%\033[38;5;253m&\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;253m&\033[38;5;250m%%\033[38;5;248m#\033[38;5;245m(\033[38;5;242m/\033[38;5;237m,\033[38;5;234m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;241m*\033[38;5;248m#\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;252m&\033[38;5;247m#\033[38;5;059m*\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;059m*\033[38;5;145m#\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;247m#\033[38;5;238m,\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;240m*\033[38;5;007m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;248m#\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;243m/\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;251m%%\033[38;5;250m%%\033[38;5;252m&\033[38;5;255m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;236m,\033[38;5;232m \033[38;5;233m \033[38;5;239m*\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m%%\033[38;5;236m,\033[38;5;232m \033[38;5;233m \033[38;5;242m/\033[38;5;254m@\033[38;5;015m@\033[38;5;254m&\033[38;5;249m%%\033[38;5;007m%%\033[38;5;253m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;007m%%\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;246m(\033[38;5;238m,\033[38;5;234m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;236m.\033[38;5;066m/\033[38;5;188m&\033[38;5;015m@\033[38;5;251m%%\033[38;5;237m,\033[38;5;232m \033[38;5;232m \033[38;5;240m*\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;249m%%\033[38;5;243m/\033[38;5;247m#\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;237m,\033[38;5;232m \033[38;5;233m \033[38;5;244m/\033[38;5;255m@\033[38;5;015m@\033[38;5;109m#\033[38;5;023m,\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;236m.\033[38;5;243m/\033[38;5;250m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;246m(\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;248m#\033[38;5;239m*\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;066m*\033[38;5;073m(\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;066m/\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;242m/\033[38;5;246m(\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;245m(\033[38;5;066m/\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;067m/\033[38;5;238m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;244m/\033[38;5;252m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m%%\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;238m,\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;240m*\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;023m*\033[38;5;074m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;074m#\033[38;5;235m.\033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;007m%%\033[38;5;250m%%\033[38;5;249m%%\033[38;5;250m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;249m%%\033[38;5;252m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;245m(\033[38;5;233m \033[38;5;016m \033[38;5;233m \033[38;5;066m*\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;236m.\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;236m.\033[38;5;245m(\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;245m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;242m/\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;023m,\033[38;5;073m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;066m*\033[38;5;233m \033[38;5;016m \033[38;5;239m*\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;244m/\033[38;5;232m \033[38;5;016m \033[38;5;235m.\033[38;5;239m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;238m,\033[38;5;236m.\033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;254m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;234m.\033[38;5;016m \033[38;5;235m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;236m,\033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;247m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;238m,\033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m,\033[38;5;016m \033[38;5;233m \033[38;5;244m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;233m \033[38;5;016m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;245m(\033[38;5;233m \033[38;5;016m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;235m.\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m*\033[38;5;232m \033[38;5;016m \033[38;5;234m.\033[38;5;246m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;238m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;243m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;241m*\033[38;5;233m \033[38;5;016m \033[38;5;237m,\033[38;5;074m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m*\033[38;5;232m \033[38;5;232m \033[38;5;244m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;145m#\033[38;5;233m \033[38;5;016m \033[38;5;239m*\033[38;5;251m%%\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;253m&\033[38;5;188m&\033[38;5;252m&\033[38;5;239m*\033[38;5;016m \033[38;5;235m.\033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;237m,\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;066m/\033[38;5;233m \033[38;5;016m \033[38;5;235m.\033[38;5;248m#\033[38;5;255m@\033[38;5;015m@\033[38;5;252m&\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;066m/\033[38;5;073m(\033[38;5;235m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;235m.\033[38;5;080m#\033[38;5;073m(\033[38;5;234m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;236m.\033[38;5;253m&\033[38;5;255m@\033[38;5;245m(\033[38;5;233m \033[38;5;016m \033[38;5;235m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;067m/\033[38;5;233m \033[38;5;232m \033[38;5;241m*\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;239m,\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;234m \033[38;5;016m \033[38;5;237m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;006m*\033[38;5;233m \033[38;5;232m \033[38;5;239m*\033[38;5;253m&\033[38;5;245m(\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;241m/\033[38;5;242m/\033[38;5;232m \033[38;5;233m \033[38;5;060m*\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;235m.\033[38;5;016m \033[38;5;236m.\033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;102m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;232m \033[38;5;233m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;235m.\033[38;5;016m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;234m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;006m*\033[38;5;232m \033[38;5;233m \033[38;5;246m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;249m#\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;238m,\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m,\033[38;5;232m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;074m#\033[38;5;235m.\033[38;5;016m \033[38;5;237m,\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;237m,\033[38;5;244m/\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;232m \033[38;5;232m \033[38;5;066m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m*\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;067m/\033[38;5;233m \033[38;5;232m \033[38;5;241m/\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m.\033[38;5;232m \033[38;5;023m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;238m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;066m/\033[38;5;233m \033[38;5;232m \033[38;5;102m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;237m,\033[38;5;016m \033[38;5;237m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;067m(\033[38;5;234m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;023m*\033[38;5;232m \033[38;5;234m.\033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;240m*\033[38;5;232m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;023m,\033[38;5;016m \033[38;5;236m.\033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;241m*\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;236m.\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;232m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;074m#\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;067m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;023m,\033[38;5;016m \033[38;5;234m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;243m/\033[38;5;232m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;067m/\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;023m*\033[38;5;232m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;253m&\033[38;5;249m%%\033[38;5;246m(\033[38;5;241m/\033[38;5;240m*\033[38;5;243m/\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;242m/\033[38;5;240m*\033[38;5;242m/\033[38;5;247m#\033[38;5;250m%%\033[38;5;188m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;242m/\033[38;5;232m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;066m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;024m*\033[38;5;232m \033[38;5;235m.\033[38;5;250m%%\033[38;5;255m@\033[38;5;252m&\033[38;5;247m#\033[38;5;242m/\033[38;5;236m.\033[38;5;234m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;234m.\033[38;5;007m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;237m,\033[38;5;243m/\033[38;5;248m#\033[38;5;253m&\033[38;5;015m@\033[38;5;254m&\033[38;5;240m*\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;060m*\033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;243m/\033[38;5;248m#\033[38;5;252m&\033[38;5;255m@\033[38;5;015m@\033[38;5;253m&\033[38;5;239m*\033[38;5;016m \033[38;5;016m \033[38;5;059m*\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;238m,\033[38;5;016m \033[38;5;232m \033[38;5;243m/\033[38;5;255m@\033[38;5;255m@\033[38;5;254m@\033[38;5;252m&\033[38;5;247m#\033[38;5;242m/\033[38;5;237m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;235m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;060m*\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;066m/\033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;239m,\033[38;5;245m(\033[38;5;251m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;234m \033[38;5;016m \033[38;5;232m \033[38;5;102m(\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;241m*\033[38;5;232m \033[38;5;016m \033[38;5;235m.\033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;250m%%\033[38;5;243m/\033[38;5;237m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;237m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;235m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;234m.\033[38;5;016m \033[38;5;242m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;242m/\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;059m*\033[38;5;253m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;007m%%\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;245m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;235m.\033[38;5;016m \033[38;5;240m*\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;067m/\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;236m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;236m,\033[38;5;016m \033[38;5;239m,\033[38;5;254m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;248m#\033[38;5;239m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;246m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;059m*\033[38;5;250m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;233m \033[38;5;232m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;067m/\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;066m*\033[38;5;232m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;241m*\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;239m*\033[38;5;250m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;247m#\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;102m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m&\033[38;5;241m*\033[38;5;232m \033[38;5;234m.\033[38;5;074m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;236m.\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;234m.\033[38;5;232m \033[38;5;243m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;252m&\033[38;5;253m&\033[38;5;255m@\033[38;5;253m&\033[38;5;246m(\033[38;5;238m,\033[38;5;236m.\033[38;5;244m(\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;243m/\033[38;5;236m.\033[38;5;239m*\033[38;5;248m#\033[38;5;254m&\033[38;5;255m@\033[38;5;252m&\033[38;5;252m&\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;250m%%\033[38;5;234m.\033[38;5;016m \033[38;5;023m*\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;023m*\033[38;5;016m \033[38;5;236m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m%%\033[38;5;239m,\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;023m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;236m.\033[38;5;243m/\033[38;5;250m%%\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;254m@\033[38;5;145m#\033[38;5;241m*\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;023m*\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;234m.\033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;238m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;249m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;247m#\033[38;5;237m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;238m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;236m.\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;233m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;236m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;251m%%\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;006m*\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;066m/\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;066m*\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;243m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;240m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;235m.\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;234m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;235m.\033[38;5;251m%%\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;234m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;067m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;235m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;067m(\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;241m*\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;188m&\033[38;5;238m,\033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m.\033[38;5;m.\033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;023m*\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;235m.\033[38;5;236m,\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;023m,\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;232m \033[38;5;235m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;m#\033[38;5;m.\033[38;5;016m \033[38;5;233m \033[38;5;248m#\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;244m/\033[38;5;232m \033[38;5;016m \033[38;5;023m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;232m \033[38;5;234m \033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;066m/\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;236m.\033[38;5;237m,\033[38;5;238m,\033[38;5;235m.\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;234m.\033[38;5;073m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;023m*\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;237m,\033[38;5;016m \033[38;5;023m,\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;073m(\033[38;5;066m/\033[38;5;066m/\033[38;5;067m/\033[38;5;073m(\033[38;5;073m(\033[38;5;234m.\033[38;5;016m \033[38;5;236m.\033[38;5;252m&\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;248m#\033[38;5;234m.\033[38;5;016m \033[38;5;234m.\033[38;5;073m(\033[38;5;074m#\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;074m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;067m/\033[38;5;233m \033[38;5;016m \033[38;5;066m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;023m*\033[38;5;074m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;067m/\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;236m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;232m \033[38;5;234m \033[38;5;067m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;235m.\033[38;5;016m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;236m.\033[38;5;238m,\033[38;5;023m*\033[38;5;238m,\033[38;5;235m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;240m*\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;195m@\033[38;5;195m@\033[38;5;159m&\033[38;5;153m&\033[38;5;153m&\033[38;5;153m&\033[38;5;153m&\033[38;5;153m&\033[38;5;195m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;252m&\033[38;5;237m,\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;235m.\033[38;5;236m.\033[38;5;237m,\033[38;5;236m,\033[38;5;235m.\033[38;5;233m \033[38;5;016m \033[38;5;232m \033[38;5;235m.\033[38;5;233m \033[38;5;016m \033[38;5;023m*\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;060m*\033[38;5;232m \033[38;5;232m \033[38;5;023m*\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;006m*\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;233m \033[38;5;066m/\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;073m(\033[38;5;235m.\033[38;5;016m \033[38;5;066m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;023m,\033[38;5;016m \033[38;5;234m \033[38;5;066m/\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;074m#\033[38;5;234m.\033[38;5;232m \033[38;5;244m/\033[38;5;255m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;255m@\033[38;5;195m&\033[38;5;117m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;153m&\033[38;5;195m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;195m@\033[38;5;195m@\033[38;5;153m&\033[38;5;153m&\033[38;5;153m&\033[38;5;159m&\033[38;5;195m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;015m@\033[38;5;253m&\033[38;5;238m,\033[38;5;016m \033[38;5;233m \033[38;5;073m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;237m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;238m,\033[38;5;016m \033[38;5;235m.\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;236m.\033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;023m,\033[38;5;073m(\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;066m/\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;236m.\033[38;5;016m \033[38;5;233m \033[38;5;102m(\033[38;5;255m@\033[38;5;195m@\033[38;5;153m&\033[38;5;117m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;153m&\033[38;5;195m&\033[38;5;195m@\033[38;5;195m@\033[38;5;195m@\033[38;5;195m@\033[38;5;195m&\033[38;5;153m&\033[38;5;117m%%\033[38;5;117m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;117m%%\033[38;5;153m&\033[38;5;195m@\033[38;5;195m@\033[38;5;195m@\033[38;5;159m&\033[38;5;153m&\033[38;5;117m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;153m&\033[38;5;159m&\033[38;5;189m&\033[38;5;159m&\033[38;5;152m&\033[38;5;066m/\033[38;5;232m \033[38;5;232m \033[38;5;023m,\033[38;5;074m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;023m*\033[38;5;066m*\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;073m(\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;236m.\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;233m \033[38;5;237m,\033[38;5;066m/\033[38;5;074m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;074m#\033[38;5;073m(\033[38;5;066m/\033[38;5;023m*\033[38;5;237m,\033[38;5;235m.\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;023m,\033[38;5;073m(\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;067m/\033[38;5;237m,\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;236m,\033[38;5;023m,\033[38;5;006m*\033[38;5;066m/\033[38;5;067m(\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;074m#\033[38;5;066m/\033[38;5;237m,\033[38;5;233m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;233m \033[38;5;236m.\033[38;5;236m.\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;234m.\033[38;5;066m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;074m(\033[38;5;023m*\033[38;5;237m,\033[38;5;023m,\033[38;5;240m*\033[38;5;066m/\033[38;5;073m(\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;067m/\033[38;5;066m/\033[38;5;060m*\033[38;5;023m*\033[38;5;060m*\033[38;5;074m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;235m.\033[38;5;235m.\033[38;5;023m,\033[38;5;023m*\033[38;5;060m*\033[38;5;023m*\033[38;5;235m.\033[38;5;232m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;232m \033[38;5;023m*\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;074m#\033[38;5;066m/\033[38;5;236m.\033[38;5;232m \033[38;5;234m.\033[38;5;067m/\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;073m(\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;074m#\033[38;5;235m.\033[38;5;232m \033[38;5;236m.\033[38;5;066m/\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;074m#\033[38;5;067m(\033[38;5;073m(\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;066m/\033[38;5;233m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;235m.\033[38;5;236m.\033[38;5;235m.\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;238m,\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;236m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;235m.\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;232m \033[38;5;016m \033[38;5;233m \033[38;5;236m.\033[38;5;066m/\033[38;5;074m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;067m/\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;067m/\033[38;5;023m,\033[38;5;234m.\033[38;5;232m \033[38;5;233m \033[38;5;234m.\033[38;5;235m.\033[38;5;238m,\033[38;5;060m*\033[38;5;066m/\033[38;5;066m/\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;073m(\033[38;5;067m/\033[38;5;066m/\033[38;5;066m/\033[38;5;023m*\033[38;5;237m,\033[38;5;235m.\033[38;5;234m.\033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;060m*\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;066m/\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;060m*\033[38;5;234m.\033[38;5;232m \033[38;5;016m \033[38;5;232m \033[38;5;234m.\033[38;5;236m.\033[38;5;023m,\033[38;5;023m*\033[38;5;066m*\033[38;5;066m*\033[38;5;066m*\033[38;5;023m,\033[38;5;237m,\033[38;5;067m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;067m/\033[38;5;237m,\033[38;5;234m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;233m \033[38;5;023m,\033[38;5;m(\033[38;5;m*\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m.\033[38;5;m(\033[38;5;m(\033[38;5;074m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;074m#\033[38;5;074m#\033[38;5;074m#\033[38;5;074m#\033[38;5;074m#\033[38;5;080m#\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;067m(\033[38;5;023m,\033[38;5;234m.\033[38;5;016m \033[38;5;233m \033[38;5;066m/\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;074m#\033[38;5;073m(\033[38;5;066m/\033[38;5;060m*\033[38;5;023m*\033[38;5;023m,\033[38;5;238m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;237m,\033[38;5;023m,\033[38;5;023m*\033[38;5;023m*\033[38;5;066m*\033[38;5;067m/\033[38;5;073m(\033[38;5;074m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m#\033[38;5;067m/\033[38;5;235m.\033[38;5;016m \033[38;5;233m \033[38;5;238m,\033[38;5;073m(\033[38;5;080m#\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;073m(\033[38;5;073m(\033[38;5;066m/\033[38;5;066m*\033[38;5;066m*\033[38;5;066m*\033[38;5;066m*\033[38;5;066m/\033[38;5;073m(\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;m%%\033[38;5;m/\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m.\033[38;5;m.\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;080m#\033[38;5;066m/\033[38;5;237m,\033[38;5;235m.\033[38;5;234m \033[38;5;233m \033[38;5;233m \033[38;5;232m \033[38;5;016m \033[38;5;016m \033[38;5;234m.\033[38;5;023m,\033[38;5;073m(\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;073m(\033[38;5;023m*\033[38;5;234m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;232m \033[38;5;233m \033[38;5;233m \033[38;5;234m \033[38;5;023m*\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;m%%\033[38;5;m#\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m.\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;m#\033[38;5;m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;081m%%\033[38;5;081m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;080m#\033[38;5;080m#\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m#\033[38;5;m*\033[38;5;m.\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m,\033[38;5;m#\033[38;5;m#\033[38;5;m%%\033[38;5;m#\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m%%\033[38;5;080m#\033[38;5;m%%\033[38;5;m%%\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m#\033[38;5;m,\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m(\033[38;5;m,\033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m \033[38;5;016m ");
	$display("\033[0");
end
endtask

endmodule
